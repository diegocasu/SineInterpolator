library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


-- ROM used to store the outputs of the SineInterpolator simulated in Python.
entity ROM_Test is
    port (
        reset : in std_logic;
        clock : in std_logic;
        address : in std_logic_vector (15 downto 0);
        data : out std_logic_vector (23 downto 0)
    );
end ROM_Test;

architecture Behaviour of ROM_Test is
 
    type rom_t is array (0 to 2**16 - 1) of std_logic_vector (23 downto 0);
    constant rom : rom_t := (
						 "000000000000000000000000",
						 "000000000000000011111111",
						 "000000000000000111111110",
						 "000000000000001011111101",
						 "000000000000001111111100",
						 "000000000000010011111011",
						 "000000000000010111111010",
						 "000000000000011011111001",
						 "000000000000011111111000",
						 "000000000000100011110111",
						 "000000000000100111110110",
						 "000000000000101011110101",
						 "000000000000101111110100",
						 "000000000000110011110011",
						 "000000000000110111110010",
						 "000000000000111011110001",
						 "000000000000000000000000",
						 "000000000000000011111111",
						 "000000000000000111111110",
						 "000000000000001011111101",
						 "000000000000001111111100",
						 "000000000000010011111011",
						 "000000000000010111111010",
						 "000000000000011011111001",
						 "000000000000011111111000",
						 "000000000000100011110111",
						 "000000000000100111110110",
						 "000000000000101011110101",
						 "000000000000101111110100",
						 "000000000000110011110011",
						 "000000000000110111110010",
						 "000000000000111011110001",
						 "000000000010100010111110",
						 "000000000010100110111101",
						 "000000000010101010111100",
						 "000000000010101110111011",
						 "000000000010110010111010",
						 "000000000010110110111001",
						 "000000000010111010111000",
						 "000000000010111110110111",
						 "000000000011000010110110",
						 "000000000011000110110101",
						 "000000000011001010110100",
						 "000000000011001110110011",
						 "000000000011010010110010",
						 "000000000011010110110001",
						 "000000000011011010110000",
						 "000000000011011110101111",
						 "000000000010100010111110",
						 "000000000010100110111101",
						 "000000000010101010111100",
						 "000000000010101110111011",
						 "000000000010110010111010",
						 "000000000010110110111001",
						 "000000000010111010111000",
						 "000000000010111110110111",
						 "000000000011000010110110",
						 "000000000011000110110101",
						 "000000000011001010110100",
						 "000000000011001110110011",
						 "000000000011010010110010",
						 "000000000011010110110001",
						 "000000000011011010110000",
						 "000000000011011110101111",
						 "000000000101000101111100",
						 "000000000101001001111011",
						 "000000000101001101111010",
						 "000000000101010001111001",
						 "000000000101010101111000",
						 "000000000101011001110111",
						 "000000000101011101110110",
						 "000000000101100001110101",
						 "000000000101100101110100",
						 "000000000101101001110011",
						 "000000000101101101110010",
						 "000000000101110001110001",
						 "000000000101110101110000",
						 "000000000101111001101111",
						 "000000000101111101101110",
						 "000000000110000001101101",
						 "000000000101000101111100",
						 "000000000101001001111011",
						 "000000000101001101111010",
						 "000000000101010001111001",
						 "000000000101010101111000",
						 "000000000101011001110111",
						 "000000000101011101110110",
						 "000000000101100001110101",
						 "000000000101100101110100",
						 "000000000101101001110011",
						 "000000000101101101110010",
						 "000000000101110001110001",
						 "000000000101110101110000",
						 "000000000101111001101111",
						 "000000000101111101101110",
						 "000000000110000001101101",
						 "000000000101000101111100",
						 "000000000101001001111011",
						 "000000000101001101111010",
						 "000000000101010001111001",
						 "000000000101010101111000",
						 "000000000101011001110111",
						 "000000000101011101110110",
						 "000000000101100001110101",
						 "000000000101100101110100",
						 "000000000101101001110011",
						 "000000000101101101110010",
						 "000000000101110001110001",
						 "000000000101110101110000",
						 "000000000101111001101111",
						 "000000000101111101101110",
						 "000000000110000001101101",
						 "000000000111101000111010",
						 "000000000111101100111001",
						 "000000000111110000111000",
						 "000000000111110100110111",
						 "000000000111111000110110",
						 "000000000111111100110101",
						 "000000001000000000110100",
						 "000000001000000100110011",
						 "000000001000001000110010",
						 "000000001000001100110001",
						 "000000001000010000110000",
						 "000000001000010100101111",
						 "000000001000011000101110",
						 "000000001000011100101101",
						 "000000001000100000101100",
						 "000000001000100100101011",
						 "000000000111101000111010",
						 "000000000111101100111001",
						 "000000000111110000111000",
						 "000000000111110100110111",
						 "000000000111111000110110",
						 "000000000111111100110101",
						 "000000001000000000110100",
						 "000000001000000100110011",
						 "000000001000001000110010",
						 "000000001000001100110001",
						 "000000001000010000110000",
						 "000000001000010100101111",
						 "000000001000011000101110",
						 "000000001000011100101101",
						 "000000001000100000101100",
						 "000000001000100100101011",
						 "000000001010001011111000",
						 "000000001010001111110111",
						 "000000001010010011110110",
						 "000000001010010111110101",
						 "000000001010011011110100",
						 "000000001010011111110011",
						 "000000001010100011110010",
						 "000000001010100111110001",
						 "000000001010101011110000",
						 "000000001010101111101111",
						 "000000001010110011101110",
						 "000000001010110111101101",
						 "000000001010111011101100",
						 "000000001010111111101011",
						 "000000001011000011101010",
						 "000000001011000111101001",
						 "000000001010001011111000",
						 "000000001010001111110111",
						 "000000001010010011110110",
						 "000000001010010111110101",
						 "000000001010011011110100",
						 "000000001010011111110011",
						 "000000001010100011110010",
						 "000000001010100111110001",
						 "000000001010101011110000",
						 "000000001010101111101111",
						 "000000001010110011101110",
						 "000000001010110111101101",
						 "000000001010111011101100",
						 "000000001010111111101011",
						 "000000001011000011101010",
						 "000000001011000111101001",
						 "000000001010001011111000",
						 "000000001010001111110111",
						 "000000001010010011110110",
						 "000000001010010111110101",
						 "000000001010011011110100",
						 "000000001010011111110011",
						 "000000001010100011110010",
						 "000000001010100111110001",
						 "000000001010101011110000",
						 "000000001010101111101111",
						 "000000001010110011101110",
						 "000000001010110111101101",
						 "000000001010111011101100",
						 "000000001010111111101011",
						 "000000001011000011101010",
						 "000000001011000111101001",
						 "000000001100101110110110",
						 "000000001100110010110101",
						 "000000001100110110110100",
						 "000000001100111010110011",
						 "000000001100111110110010",
						 "000000001101000010110001",
						 "000000001101000110110000",
						 "000000001101001010101111",
						 "000000001101001110101110",
						 "000000001101010010101101",
						 "000000001101010110101100",
						 "000000001101011010101011",
						 "000000001101011110101010",
						 "000000001101100010101001",
						 "000000001101100110101000",
						 "000000001101101010100111",
						 "000000001100101110110110",
						 "000000001100110010110101",
						 "000000001100110110110100",
						 "000000001100111010110011",
						 "000000001100111110110010",
						 "000000001101000010110001",
						 "000000001101000110110000",
						 "000000001101001010101111",
						 "000000001101001110101110",
						 "000000001101010010101101",
						 "000000001101010110101100",
						 "000000001101011010101011",
						 "000000001101011110101010",
						 "000000001101100010101001",
						 "000000001101100110101000",
						 "000000001101101010100111",
						 "000000001100101110110110",
						 "000000001100110010110101",
						 "000000001100110110110100",
						 "000000001100111010110011",
						 "000000001100111110110010",
						 "000000001101000010110001",
						 "000000001101000110110000",
						 "000000001101001010101111",
						 "000000001101001110101110",
						 "000000001101010010101101",
						 "000000001101010110101100",
						 "000000001101011010101011",
						 "000000001101011110101010",
						 "000000001101100010101001",
						 "000000001101100110101000",
						 "000000001101101010100111",
						 "000000001111010001110100",
						 "000000001111010101110011",
						 "000000001111011001110010",
						 "000000001111011101110001",
						 "000000001111100001110000",
						 "000000001111100101101111",
						 "000000001111101001101110",
						 "000000001111101101101101",
						 "000000001111110001101100",
						 "000000001111110101101011",
						 "000000001111111001101010",
						 "000000001111111101101001",
						 "000000010000000001101000",
						 "000000010000000101100111",
						 "000000010000001001100110",
						 "000000010000001101100101",
						 "000000001111010001110100",
						 "000000001111010101110011",
						 "000000001111011001110010",
						 "000000001111011101110001",
						 "000000001111100001110000",
						 "000000001111100101101111",
						 "000000001111101001101110",
						 "000000001111101101101101",
						 "000000001111110001101100",
						 "000000001111110101101011",
						 "000000001111111001101010",
						 "000000001111111101101001",
						 "000000010000000001101000",
						 "000000010000000101100111",
						 "000000010000001001100110",
						 "000000010000001101100101",
						 "000000010001110100110010",
						 "000000010001111000110001",
						 "000000010001111100110000",
						 "000000010010000000101111",
						 "000000010010000100101110",
						 "000000010010001000101101",
						 "000000010010001100101100",
						 "000000010010010000101011",
						 "000000010010010100101010",
						 "000000010010011000101001",
						 "000000010010011100101000",
						 "000000010010100000100111",
						 "000000010010100100100110",
						 "000000010010101000100101",
						 "000000010010101100100100",
						 "000000010010110000100011",
						 "000000010001110100110010",
						 "000000010001111000110001",
						 "000000010001111100110000",
						 "000000010010000000101111",
						 "000000010010000100101110",
						 "000000010010001000101101",
						 "000000010010001100101100",
						 "000000010010010000101011",
						 "000000010010010100101010",
						 "000000010010011000101001",
						 "000000010010011100101000",
						 "000000010010100000100111",
						 "000000010010100100100110",
						 "000000010010101000100101",
						 "000000010010101100100100",
						 "000000010010110000100011",
						 "000000010001110100110010",
						 "000000010001111000110001",
						 "000000010001111100110000",
						 "000000010010000000101111",
						 "000000010010000100101110",
						 "000000010010001000101101",
						 "000000010010001100101100",
						 "000000010010010000101011",
						 "000000010010010100101010",
						 "000000010010011000101001",
						 "000000010010011100101000",
						 "000000010010100000100111",
						 "000000010010100100100110",
						 "000000010010101000100101",
						 "000000010010101100100100",
						 "000000010010110000100011",
						 "000000010100010111110000",
						 "000000010100011011101111",
						 "000000010100011111101110",
						 "000000010100100011101101",
						 "000000010100100111101100",
						 "000000010100101011101011",
						 "000000010100101111101010",
						 "000000010100110011101001",
						 "000000010100110111101000",
						 "000000010100111011100111",
						 "000000010100111111100110",
						 "000000010101000011100101",
						 "000000010101000111100100",
						 "000000010101001011100011",
						 "000000010101001111100010",
						 "000000010101010011100001",
						 "000000010100010111110000",
						 "000000010100011011101111",
						 "000000010100011111101110",
						 "000000010100100011101101",
						 "000000010100100111101100",
						 "000000010100101011101011",
						 "000000010100101111101010",
						 "000000010100110011101001",
						 "000000010100110111101000",
						 "000000010100111011100111",
						 "000000010100111111100110",
						 "000000010101000011100101",
						 "000000010101000111100100",
						 "000000010101001011100011",
						 "000000010101001111100010",
						 "000000010101010011100001",
						 "000000010110111010101110",
						 "000000010110111110101101",
						 "000000010111000010101100",
						 "000000010111000110101011",
						 "000000010111001010101010",
						 "000000010111001110101001",
						 "000000010111010010101000",
						 "000000010111010110100111",
						 "000000010111011010100110",
						 "000000010111011110100101",
						 "000000010111100010100100",
						 "000000010111100110100011",
						 "000000010111101010100010",
						 "000000010111101110100001",
						 "000000010111110010100000",
						 "000000010111110110011111",
						 "000000010110111010101110",
						 "000000010110111110101101",
						 "000000010111000010101100",
						 "000000010111000110101011",
						 "000000010111001010101010",
						 "000000010111001110101001",
						 "000000010111010010101000",
						 "000000010111010110100111",
						 "000000010111011010100110",
						 "000000010111011110100101",
						 "000000010111100010100100",
						 "000000010111100110100011",
						 "000000010111101010100010",
						 "000000010111101110100001",
						 "000000010111110010100000",
						 "000000010111110110011111",
						 "000000010110111010101110",
						 "000000010110111110101101",
						 "000000010111000010101100",
						 "000000010111000110101011",
						 "000000010111001010101010",
						 "000000010111001110101001",
						 "000000010111010010101000",
						 "000000010111010110100111",
						 "000000010111011010100110",
						 "000000010111011110100101",
						 "000000010111100010100100",
						 "000000010111100110100011",
						 "000000010111101010100010",
						 "000000010111101110100001",
						 "000000010111110010100000",
						 "000000010111110110011111",
						 "000000011001011101101100",
						 "000000011001100001101011",
						 "000000011001100101101010",
						 "000000011001101001101001",
						 "000000011001101101101000",
						 "000000011001110001100111",
						 "000000011001110101100110",
						 "000000011001111001100101",
						 "000000011001111101100100",
						 "000000011010000001100011",
						 "000000011010000101100010",
						 "000000011010001001100001",
						 "000000011010001101100000",
						 "000000011010010001011111",
						 "000000011010010101011110",
						 "000000011010011001011101",
						 "000000011001011101101100",
						 "000000011001100001101011",
						 "000000011001100101101010",
						 "000000011001101001101001",
						 "000000011001101101101000",
						 "000000011001110001100111",
						 "000000011001110101100110",
						 "000000011001111001100101",
						 "000000011001111101100100",
						 "000000011010000001100011",
						 "000000011010000101100010",
						 "000000011010001001100001",
						 "000000011010001101100000",
						 "000000011010010001011111",
						 "000000011010010101011110",
						 "000000011010011001011101",
						 "000000011100000000101010",
						 "000000011100000100101001",
						 "000000011100001000101000",
						 "000000011100001100100111",
						 "000000011100010000100110",
						 "000000011100010100100101",
						 "000000011100011000100100",
						 "000000011100011100100011",
						 "000000011100100000100010",
						 "000000011100100100100001",
						 "000000011100101000100000",
						 "000000011100101100011111",
						 "000000011100110000011110",
						 "000000011100110100011101",
						 "000000011100111000011100",
						 "000000011100111100011011",
						 "000000011100000000101010",
						 "000000011100000100101001",
						 "000000011100001000101000",
						 "000000011100001100100111",
						 "000000011100010000100110",
						 "000000011100010100100101",
						 "000000011100011000100100",
						 "000000011100011100100011",
						 "000000011100100000100010",
						 "000000011100100100100001",
						 "000000011100101000100000",
						 "000000011100101100011111",
						 "000000011100110000011110",
						 "000000011100110100011101",
						 "000000011100111000011100",
						 "000000011100111100011011",
						 "000000011100000000101010",
						 "000000011100000100101001",
						 "000000011100001000101000",
						 "000000011100001100100111",
						 "000000011100010000100110",
						 "000000011100010100100101",
						 "000000011100011000100100",
						 "000000011100011100100011",
						 "000000011100100000100010",
						 "000000011100100100100001",
						 "000000011100101000100000",
						 "000000011100101100011111",
						 "000000011100110000011110",
						 "000000011100110100011101",
						 "000000011100111000011100",
						 "000000011100111100011011",
						 "000000011110100011101000",
						 "000000011110100111100111",
						 "000000011110101011100110",
						 "000000011110101111100101",
						 "000000011110110011100100",
						 "000000011110110111100011",
						 "000000011110111011100010",
						 "000000011110111111100001",
						 "000000011111000011100000",
						 "000000011111000111011111",
						 "000000011111001011011110",
						 "000000011111001111011101",
						 "000000011111010011011100",
						 "000000011111010111011011",
						 "000000011111011011011010",
						 "000000011111011111011001",
						 "000000011110100011101000",
						 "000000011110100111100111",
						 "000000011110101011100110",
						 "000000011110101111100101",
						 "000000011110110011100100",
						 "000000011110110111100011",
						 "000000011110111011100010",
						 "000000011110111111100001",
						 "000000011111000011100000",
						 "000000011111000111011111",
						 "000000011111001011011110",
						 "000000011111001111011101",
						 "000000011111010011011100",
						 "000000011111010111011011",
						 "000000011111011011011010",
						 "000000011111011111011001",
						 "000000100001000110100110",
						 "000000100001001010100101",
						 "000000100001001110100100",
						 "000000100001010010100011",
						 "000000100001010110100010",
						 "000000100001011010100001",
						 "000000100001011110100000",
						 "000000100001100010011111",
						 "000000100001100110011110",
						 "000000100001101010011101",
						 "000000100001101110011100",
						 "000000100001110010011011",
						 "000000100001110110011010",
						 "000000100001111010011001",
						 "000000100001111110011000",
						 "000000100010000010010111",
						 "000000100001000110100110",
						 "000000100001001010100101",
						 "000000100001001110100100",
						 "000000100001010010100011",
						 "000000100001010110100010",
						 "000000100001011010100001",
						 "000000100001011110100000",
						 "000000100001100010011111",
						 "000000100001100110011110",
						 "000000100001101010011101",
						 "000000100001101110011100",
						 "000000100001110010011011",
						 "000000100001110110011010",
						 "000000100001111010011001",
						 "000000100001111110011000",
						 "000000100010000010010111",
						 "000000100001000110100110",
						 "000000100001001010100101",
						 "000000100001001110100100",
						 "000000100001010010100011",
						 "000000100001010110100010",
						 "000000100001011010100001",
						 "000000100001011110100000",
						 "000000100001100010011111",
						 "000000100001100110011110",
						 "000000100001101010011101",
						 "000000100001101110011100",
						 "000000100001110010011011",
						 "000000100001110110011010",
						 "000000100001111010011001",
						 "000000100001111110011000",
						 "000000100010000010010111",
						 "000000100011101001100100",
						 "000000100011101101100011",
						 "000000100011110001100010",
						 "000000100011110101100001",
						 "000000100011111001100000",
						 "000000100011111101011111",
						 "000000100100000001011110",
						 "000000100100000101011101",
						 "000000100100001001011100",
						 "000000100100001101011011",
						 "000000100100010001011010",
						 "000000100100010101011001",
						 "000000100100011001011000",
						 "000000100100011101010111",
						 "000000100100100001010110",
						 "000000100100100101010101",
						 "000000100011101001100100",
						 "000000100011101101100011",
						 "000000100011110001100010",
						 "000000100011110101100001",
						 "000000100011111001100000",
						 "000000100011111101011111",
						 "000000100100000001011110",
						 "000000100100000101011101",
						 "000000100100001001011100",
						 "000000100100001101011011",
						 "000000100100010001011010",
						 "000000100100010101011001",
						 "000000100100011001011000",
						 "000000100100011101010111",
						 "000000100100100001010110",
						 "000000100100100101010101",
						 "000000100011101001100100",
						 "000000100011101101100011",
						 "000000100011110001100010",
						 "000000100011110101100001",
						 "000000100011111001100000",
						 "000000100011111101011111",
						 "000000100100000001011110",
						 "000000100100000101011101",
						 "000000100100001001011100",
						 "000000100100001101011011",
						 "000000100100010001011010",
						 "000000100100010101011001",
						 "000000100100011001011000",
						 "000000100100011101010111",
						 "000000100100100001010110",
						 "000000100100100101010101",
						 "000000100110001100100010",
						 "000000100110010000100001",
						 "000000100110010100100000",
						 "000000100110011000011111",
						 "000000100110011100011110",
						 "000000100110100000011101",
						 "000000100110100100011100",
						 "000000100110101000011011",
						 "000000100110101100011010",
						 "000000100110110000011001",
						 "000000100110110100011000",
						 "000000100110111000010111",
						 "000000100110111100010110",
						 "000000100111000000010101",
						 "000000100111000100010100",
						 "000000100111001000010011",
						 "000000100110001100100010",
						 "000000100110010000100001",
						 "000000100110010100100000",
						 "000000100110011000011111",
						 "000000100110011100011110",
						 "000000100110100000011101",
						 "000000100110100100011100",
						 "000000100110101000011011",
						 "000000100110101100011010",
						 "000000100110110000011001",
						 "000000100110110100011000",
						 "000000100110111000010111",
						 "000000100110111100010110",
						 "000000100111000000010101",
						 "000000100111000100010100",
						 "000000100111001000010011",
						 "000000101000101111100000",
						 "000000101000110011011111",
						 "000000101000110111011110",
						 "000000101000111011011101",
						 "000000101000111111011100",
						 "000000101001000011011011",
						 "000000101001000111011010",
						 "000000101001001011011001",
						 "000000101001001111011000",
						 "000000101001010011010111",
						 "000000101001010111010110",
						 "000000101001011011010101",
						 "000000101001011111010100",
						 "000000101001100011010011",
						 "000000101001100111010010",
						 "000000101001101011010001",
						 "000000101000101111100000",
						 "000000101000110011011110",
						 "000000101000110111011100",
						 "000000101000111011011010",
						 "000000101000111111011000",
						 "000000101001000011010110",
						 "000000101001000111010100",
						 "000000101001001011010010",
						 "000000101001001111010000",
						 "000000101001010011001110",
						 "000000101001010111001100",
						 "000000101001011011001010",
						 "000000101001011111001000",
						 "000000101001100011000110",
						 "000000101001100111000100",
						 "000000101001101011000010",
						 "000000101000101111100000",
						 "000000101000110011011110",
						 "000000101000110111011100",
						 "000000101000111011011010",
						 "000000101000111111011000",
						 "000000101001000011010110",
						 "000000101001000111010100",
						 "000000101001001011010010",
						 "000000101001001111010000",
						 "000000101001010011001110",
						 "000000101001010111001100",
						 "000000101001011011001010",
						 "000000101001011111001000",
						 "000000101001100011000110",
						 "000000101001100111000100",
						 "000000101001101011000010",
						 "000000101011010010011110",
						 "000000101011010110011100",
						 "000000101011011010011010",
						 "000000101011011110011000",
						 "000000101011100010010110",
						 "000000101011100110010100",
						 "000000101011101010010010",
						 "000000101011101110010000",
						 "000000101011110010001110",
						 "000000101011110110001100",
						 "000000101011111010001010",
						 "000000101011111110001000",
						 "000000101100000010000110",
						 "000000101100000110000100",
						 "000000101100001010000010",
						 "000000101100001110000000",
						 "000000101011010010011110",
						 "000000101011010110011100",
						 "000000101011011010011010",
						 "000000101011011110011000",
						 "000000101011100010010110",
						 "000000101011100110010100",
						 "000000101011101010010010",
						 "000000101011101110010000",
						 "000000101011110010001110",
						 "000000101011110110001100",
						 "000000101011111010001010",
						 "000000101011111110001000",
						 "000000101100000010000110",
						 "000000101100000110000100",
						 "000000101100001010000010",
						 "000000101100001110000000",
						 "000000101101110101011100",
						 "000000101101111001011010",
						 "000000101101111101011000",
						 "000000101110000001010110",
						 "000000101110000101010100",
						 "000000101110001001010010",
						 "000000101110001101010000",
						 "000000101110010001001110",
						 "000000101110010101001100",
						 "000000101110011001001010",
						 "000000101110011101001000",
						 "000000101110100001000110",
						 "000000101110100101000100",
						 "000000101110101001000010",
						 "000000101110101101000000",
						 "000000101110110000111110",
						 "000000101101110101011100",
						 "000000101101111001011010",
						 "000000101101111101011000",
						 "000000101110000001010110",
						 "000000101110000101010100",
						 "000000101110001001010010",
						 "000000101110001101010000",
						 "000000101110010001001110",
						 "000000101110010101001100",
						 "000000101110011001001010",
						 "000000101110011101001000",
						 "000000101110100001000110",
						 "000000101110100101000100",
						 "000000101110101001000010",
						 "000000101110101101000000",
						 "000000101110110000111110",
						 "000000101101110101011100",
						 "000000101101111001011010",
						 "000000101101111101011000",
						 "000000101110000001010110",
						 "000000101110000101010100",
						 "000000101110001001010010",
						 "000000101110001101010000",
						 "000000101110010001001110",
						 "000000101110010101001100",
						 "000000101110011001001010",
						 "000000101110011101001000",
						 "000000101110100001000110",
						 "000000101110100101000100",
						 "000000101110101001000010",
						 "000000101110101101000000",
						 "000000101110110000111110",
						 "000000110000011000011010",
						 "000000110000011100011000",
						 "000000110000100000010110",
						 "000000110000100100010100",
						 "000000110000101000010010",
						 "000000110000101100010000",
						 "000000110000110000001110",
						 "000000110000110100001100",
						 "000000110000111000001010",
						 "000000110000111100001000",
						 "000000110001000000000110",
						 "000000110001000100000100",
						 "000000110001001000000010",
						 "000000110001001100000000",
						 "000000110001001111111110",
						 "000000110001010011111100",
						 "000000110000011000011010",
						 "000000110000011100011000",
						 "000000110000100000010110",
						 "000000110000100100010100",
						 "000000110000101000010010",
						 "000000110000101100010000",
						 "000000110000110000001110",
						 "000000110000110100001100",
						 "000000110000111000001010",
						 "000000110000111100001000",
						 "000000110001000000000110",
						 "000000110001000100000100",
						 "000000110001001000000010",
						 "000000110001001100000000",
						 "000000110001001111111110",
						 "000000110001010011111100",
						 "000000110010111011011000",
						 "000000110010111111010110",
						 "000000110011000011010100",
						 "000000110011000111010010",
						 "000000110011001011010000",
						 "000000110011001111001110",
						 "000000110011010011001100",
						 "000000110011010111001010",
						 "000000110011011011001000",
						 "000000110011011111000110",
						 "000000110011100011000100",
						 "000000110011100111000010",
						 "000000110011101011000000",
						 "000000110011101110111110",
						 "000000110011110010111100",
						 "000000110011110110111010",
						 "000000110010111011011000",
						 "000000110010111111010110",
						 "000000110011000011010100",
						 "000000110011000111010010",
						 "000000110011001011010000",
						 "000000110011001111001110",
						 "000000110011010011001100",
						 "000000110011010111001010",
						 "000000110011011011001000",
						 "000000110011011111000110",
						 "000000110011100011000100",
						 "000000110011100111000010",
						 "000000110011101011000000",
						 "000000110011101110111110",
						 "000000110011110010111100",
						 "000000110011110110111010",
						 "000000110010111011011000",
						 "000000110010111111010110",
						 "000000110011000011010100",
						 "000000110011000111010010",
						 "000000110011001011010000",
						 "000000110011001111001110",
						 "000000110011010011001100",
						 "000000110011010111001010",
						 "000000110011011011001000",
						 "000000110011011111000110",
						 "000000110011100011000100",
						 "000000110011100111000010",
						 "000000110011101011000000",
						 "000000110011101110111110",
						 "000000110011110010111100",
						 "000000110011110110111010",
						 "000000110101011110010110",
						 "000000110101100010010100",
						 "000000110101100110010010",
						 "000000110101101010010000",
						 "000000110101101110001110",
						 "000000110101110010001100",
						 "000000110101110110001010",
						 "000000110101111010001000",
						 "000000110101111110000110",
						 "000000110110000010000100",
						 "000000110110000110000010",
						 "000000110110001010000000",
						 "000000110110001101111110",
						 "000000110110010001111100",
						 "000000110110010101111010",
						 "000000110110011001111000",
						 "000000110101011110010110",
						 "000000110101100010010100",
						 "000000110101100110010010",
						 "000000110101101010010000",
						 "000000110101101110001110",
						 "000000110101110010001100",
						 "000000110101110110001010",
						 "000000110101111010001000",
						 "000000110101111110000110",
						 "000000110110000010000100",
						 "000000110110000110000010",
						 "000000110110001010000000",
						 "000000110110001101111110",
						 "000000110110010001111100",
						 "000000110110010101111010",
						 "000000110110011001111000",
						 "000000110101011110010110",
						 "000000110101100010010100",
						 "000000110101100110010010",
						 "000000110101101010010000",
						 "000000110101101110001110",
						 "000000110101110010001100",
						 "000000110101110110001010",
						 "000000110101111010001000",
						 "000000110101111110000110",
						 "000000110110000010000100",
						 "000000110110000110000010",
						 "000000110110001010000000",
						 "000000110110001101111110",
						 "000000110110010001111100",
						 "000000110110010101111010",
						 "000000110110011001111000",
						 "000000111000000001010100",
						 "000000111000000101010010",
						 "000000111000001001010000",
						 "000000111000001101001110",
						 "000000111000010001001100",
						 "000000111000010101001010",
						 "000000111000011001001000",
						 "000000111000011101000110",
						 "000000111000100001000100",
						 "000000111000100101000010",
						 "000000111000101001000000",
						 "000000111000101100111110",
						 "000000111000110000111100",
						 "000000111000110100111010",
						 "000000111000111000111000",
						 "000000111000111100110110",
						 "000000111000000001010100",
						 "000000111000000101010010",
						 "000000111000001001010000",
						 "000000111000001101001110",
						 "000000111000010001001100",
						 "000000111000010101001010",
						 "000000111000011001001000",
						 "000000111000011101000110",
						 "000000111000100001000100",
						 "000000111000100101000010",
						 "000000111000101001000000",
						 "000000111000101100111110",
						 "000000111000110000111100",
						 "000000111000110100111010",
						 "000000111000111000111000",
						 "000000111000111100110110",
						 "000000111010100100010010",
						 "000000111010101000010000",
						 "000000111010101100001110",
						 "000000111010110000001100",
						 "000000111010110100001010",
						 "000000111010111000001000",
						 "000000111010111100000110",
						 "000000111011000000000100",
						 "000000111011000100000010",
						 "000000111011001000000000",
						 "000000111011001011111110",
						 "000000111011001111111100",
						 "000000111011010011111010",
						 "000000111011010111111000",
						 "000000111011011011110110",
						 "000000111011011111110100",
						 "000000111010100100010010",
						 "000000111010101000010000",
						 "000000111010101100001110",
						 "000000111010110000001100",
						 "000000111010110100001010",
						 "000000111010111000001000",
						 "000000111010111100000110",
						 "000000111011000000000100",
						 "000000111011000100000010",
						 "000000111011001000000000",
						 "000000111011001011111110",
						 "000000111011001111111100",
						 "000000111011010011111010",
						 "000000111011010111111000",
						 "000000111011011011110110",
						 "000000111011011111110100",
						 "000000111010100100010010",
						 "000000111010101000010000",
						 "000000111010101100001110",
						 "000000111010110000001100",
						 "000000111010110100001010",
						 "000000111010111000001000",
						 "000000111010111100000110",
						 "000000111011000000000100",
						 "000000111011000100000010",
						 "000000111011001000000000",
						 "000000111011001011111110",
						 "000000111011001111111100",
						 "000000111011010011111010",
						 "000000111011010111111000",
						 "000000111011011011110110",
						 "000000111011011111110100",
						 "000000111101000111010000",
						 "000000111101001011001110",
						 "000000111101001111001100",
						 "000000111101010011001010",
						 "000000111101010111001000",
						 "000000111101011011000110",
						 "000000111101011111000100",
						 "000000111101100011000010",
						 "000000111101100111000000",
						 "000000111101101010111110",
						 "000000111101101110111100",
						 "000000111101110010111010",
						 "000000111101110110111000",
						 "000000111101111010110110",
						 "000000111101111110110100",
						 "000000111110000010110010",
						 "000000111101000111010000",
						 "000000111101001011001110",
						 "000000111101001111001100",
						 "000000111101010011001010",
						 "000000111101010111001000",
						 "000000111101011011000110",
						 "000000111101011111000100",
						 "000000111101100011000010",
						 "000000111101100111000000",
						 "000000111101101010111110",
						 "000000111101101110111100",
						 "000000111101110010111010",
						 "000000111101110110111000",
						 "000000111101111010110110",
						 "000000111101111110110100",
						 "000000111110000010110010",
						 "000000111111101010001110",
						 "000000111111101110001100",
						 "000000111111110010001010",
						 "000000111111110110001000",
						 "000000111111111010000110",
						 "000000111111111110000100",
						 "000001000000000010000010",
						 "000001000000000110000000",
						 "000001000000001001111110",
						 "000001000000001101111100",
						 "000001000000010001111010",
						 "000001000000010101111000",
						 "000001000000011001110110",
						 "000001000000011101110100",
						 "000001000000100001110010",
						 "000001000000100101110000",
						 "000000111111101010001110",
						 "000000111111101110001100",
						 "000000111111110010001010",
						 "000000111111110110001000",
						 "000000111111111010000110",
						 "000000111111111110000100",
						 "000001000000000010000010",
						 "000001000000000110000000",
						 "000001000000001001111110",
						 "000001000000001101111100",
						 "000001000000010001111010",
						 "000001000000010101111000",
						 "000001000000011001110110",
						 "000001000000011101110100",
						 "000001000000100001110010",
						 "000001000000100101110000",
						 "000000111111101010001110",
						 "000000111111101110001100",
						 "000000111111110010001010",
						 "000000111111110110001000",
						 "000000111111111010000110",
						 "000000111111111110000100",
						 "000001000000000010000010",
						 "000001000000000110000000",
						 "000001000000001001111110",
						 "000001000000001101111100",
						 "000001000000010001111010",
						 "000001000000010101111000",
						 "000001000000011001110110",
						 "000001000000011101110100",
						 "000001000000100001110010",
						 "000001000000100101110000",
						 "000001000010001101001100",
						 "000001000010010001001010",
						 "000001000010010101001000",
						 "000001000010011001000110",
						 "000001000010011101000100",
						 "000001000010100001000010",
						 "000001000010100101000000",
						 "000001000010101000111110",
						 "000001000010101100111100",
						 "000001000010110000111010",
						 "000001000010110100111000",
						 "000001000010111000110110",
						 "000001000010111100110100",
						 "000001000011000000110010",
						 "000001000011000100110000",
						 "000001000011001000101110",
						 "000001000010001101001100",
						 "000001000010010001001010",
						 "000001000010010101001000",
						 "000001000010011001000110",
						 "000001000010011101000100",
						 "000001000010100001000010",
						 "000001000010100101000000",
						 "000001000010101000111110",
						 "000001000010101100111100",
						 "000001000010110000111010",
						 "000001000010110100111000",
						 "000001000010111000110110",
						 "000001000010111100110100",
						 "000001000011000000110010",
						 "000001000011000100110000",
						 "000001000011001000101110",
						 "000001000100110000001010",
						 "000001000100110100001000",
						 "000001000100111000000110",
						 "000001000100111100000100",
						 "000001000101000000000010",
						 "000001000101000100000000",
						 "000001000101000111111110",
						 "000001000101001011111100",
						 "000001000101001111111010",
						 "000001000101010011111000",
						 "000001000101010111110110",
						 "000001000101011011110100",
						 "000001000101011111110010",
						 "000001000101100011110000",
						 "000001000101100111101110",
						 "000001000101101011101100",
						 "000001000100110000001010",
						 "000001000100110100001000",
						 "000001000100111000000110",
						 "000001000100111100000100",
						 "000001000101000000000010",
						 "000001000101000100000000",
						 "000001000101000111111110",
						 "000001000101001011111100",
						 "000001000101001111111010",
						 "000001000101010011111000",
						 "000001000101010111110110",
						 "000001000101011011110100",
						 "000001000101011111110010",
						 "000001000101100011110000",
						 "000001000101100111101110",
						 "000001000101101011101100",
						 "000001000100110000001010",
						 "000001000100110100001000",
						 "000001000100111000000110",
						 "000001000100111100000100",
						 "000001000101000000000010",
						 "000001000101000100000000",
						 "000001000101000111111110",
						 "000001000101001011111100",
						 "000001000101001111111010",
						 "000001000101010011111000",
						 "000001000101010111110110",
						 "000001000101011011110100",
						 "000001000101011111110010",
						 "000001000101100011110000",
						 "000001000101100111101110",
						 "000001000101101011101100",
						 "000001000111010011001000",
						 "000001000111010111000101",
						 "000001000111011011000010",
						 "000001000111011110111111",
						 "000001000111100010111100",
						 "000001000111100110111001",
						 "000001000111101010110110",
						 "000001000111101110110011",
						 "000001000111110010110000",
						 "000001000111110110101101",
						 "000001000111111010101010",
						 "000001000111111110100111",
						 "000001001000000010100100",
						 "000001001000000110100001",
						 "000001001000001010011110",
						 "000001001000001110011011",
						 "000001000111010011001000",
						 "000001000111010111000101",
						 "000001000111011011000010",
						 "000001000111011110111111",
						 "000001000111100010111100",
						 "000001000111100110111001",
						 "000001000111101010110110",
						 "000001000111101110110011",
						 "000001000111110010110000",
						 "000001000111110110101101",
						 "000001000111111010101010",
						 "000001000111111110100111",
						 "000001001000000010100100",
						 "000001001000000110100001",
						 "000001001000001010011110",
						 "000001001000001110011011",
						 "000001000111010011001000",
						 "000001000111010111000101",
						 "000001000111011011000010",
						 "000001000111011110111111",
						 "000001000111100010111100",
						 "000001000111100110111001",
						 "000001000111101010110110",
						 "000001000111101110110011",
						 "000001000111110010110000",
						 "000001000111110110101101",
						 "000001000111111010101010",
						 "000001000111111110100111",
						 "000001001000000010100100",
						 "000001001000000110100001",
						 "000001001000001010011110",
						 "000001001000001110011011",
						 "000001001001110110000110",
						 "000001001001111010000011",
						 "000001001001111110000000",
						 "000001001010000001111101",
						 "000001001010000101111010",
						 "000001001010001001110111",
						 "000001001010001101110100",
						 "000001001010010001110001",
						 "000001001010010101101110",
						 "000001001010011001101011",
						 "000001001010011101101000",
						 "000001001010100001100101",
						 "000001001010100101100010",
						 "000001001010101001011111",
						 "000001001010101101011100",
						 "000001001010110001011001",
						 "000001001001110110000110",
						 "000001001001111010000011",
						 "000001001001111110000000",
						 "000001001010000001111101",
						 "000001001010000101111010",
						 "000001001010001001110111",
						 "000001001010001101110100",
						 "000001001010010001110001",
						 "000001001010010101101110",
						 "000001001010011001101011",
						 "000001001010011101101000",
						 "000001001010100001100101",
						 "000001001010100101100010",
						 "000001001010101001011111",
						 "000001001010101101011100",
						 "000001001010110001011001",
						 "000001001100011001000100",
						 "000001001100011101000001",
						 "000001001100100000111110",
						 "000001001100100100111011",
						 "000001001100101000111000",
						 "000001001100101100110101",
						 "000001001100110000110010",
						 "000001001100110100101111",
						 "000001001100111000101100",
						 "000001001100111100101001",
						 "000001001101000000100110",
						 "000001001101000100100011",
						 "000001001101001000100000",
						 "000001001101001100011101",
						 "000001001101010000011010",
						 "000001001101010100010111",
						 "000001001100011001000100",
						 "000001001100011101000001",
						 "000001001100100000111110",
						 "000001001100100100111011",
						 "000001001100101000111000",
						 "000001001100101100110101",
						 "000001001100110000110010",
						 "000001001100110100101111",
						 "000001001100111000101100",
						 "000001001100111100101001",
						 "000001001101000000100110",
						 "000001001101000100100011",
						 "000001001101001000100000",
						 "000001001101001100011101",
						 "000001001101010000011010",
						 "000001001101010100010111",
						 "000001001100011001000100",
						 "000001001100011101000001",
						 "000001001100100000111110",
						 "000001001100100100111011",
						 "000001001100101000111000",
						 "000001001100101100110101",
						 "000001001100110000110010",
						 "000001001100110100101111",
						 "000001001100111000101100",
						 "000001001100111100101001",
						 "000001001101000000100110",
						 "000001001101000100100011",
						 "000001001101001000100000",
						 "000001001101001100011101",
						 "000001001101010000011010",
						 "000001001101010100010111",
						 "000001001110111100000010",
						 "000001001110111111111111",
						 "000001001111000011111100",
						 "000001001111000111111001",
						 "000001001111001011110110",
						 "000001001111001111110011",
						 "000001001111010011110000",
						 "000001001111010111101101",
						 "000001001111011011101010",
						 "000001001111011111100111",
						 "000001001111100011100100",
						 "000001001111100111100001",
						 "000001001111101011011110",
						 "000001001111101111011011",
						 "000001001111110011011000",
						 "000001001111110111010101",
						 "000001001110111100000010",
						 "000001001110111111111111",
						 "000001001111000011111100",
						 "000001001111000111111001",
						 "000001001111001011110110",
						 "000001001111001111110011",
						 "000001001111010011110000",
						 "000001001111010111101101",
						 "000001001111011011101010",
						 "000001001111011111100111",
						 "000001001111100011100100",
						 "000001001111100111100001",
						 "000001001111101011011110",
						 "000001001111101111011011",
						 "000001001111110011011000",
						 "000001001111110111010101",
						 "000001010001011111000000",
						 "000001010001100010111101",
						 "000001010001100110111010",
						 "000001010001101010110111",
						 "000001010001101110110100",
						 "000001010001110010110001",
						 "000001010001110110101110",
						 "000001010001111010101011",
						 "000001010001111110101000",
						 "000001010010000010100101",
						 "000001010010000110100010",
						 "000001010010001010011111",
						 "000001010010001110011100",
						 "000001010010010010011001",
						 "000001010010010110010110",
						 "000001010010011010010011",
						 "000001010001011111000000",
						 "000001010001100010111101",
						 "000001010001100110111010",
						 "000001010001101010110111",
						 "000001010001101110110100",
						 "000001010001110010110001",
						 "000001010001110110101110",
						 "000001010001111010101011",
						 "000001010001111110101000",
						 "000001010010000010100101",
						 "000001010010000110100010",
						 "000001010010001010011111",
						 "000001010010001110011100",
						 "000001010010010010011001",
						 "000001010010010110010110",
						 "000001010010011010010011",
						 "000001010001011111000000",
						 "000001010001100010111101",
						 "000001010001100110111010",
						 "000001010001101010110111",
						 "000001010001101110110100",
						 "000001010001110010110001",
						 "000001010001110110101110",
						 "000001010001111010101011",
						 "000001010001111110101000",
						 "000001010010000010100101",
						 "000001010010000110100010",
						 "000001010010001010011111",
						 "000001010010001110011100",
						 "000001010010010010011001",
						 "000001010010010110010110",
						 "000001010010011010010011",
						 "000001010100000001111110",
						 "000001010100000101111011",
						 "000001010100001001111000",
						 "000001010100001101110101",
						 "000001010100010001110010",
						 "000001010100010101101111",
						 "000001010100011001101100",
						 "000001010100011101101001",
						 "000001010100100001100110",
						 "000001010100100101100011",
						 "000001010100101001100000",
						 "000001010100101101011101",
						 "000001010100110001011010",
						 "000001010100110101010111",
						 "000001010100111001010100",
						 "000001010100111101010001",
						 "000001010100000001111110",
						 "000001010100000101111011",
						 "000001010100001001111000",
						 "000001010100001101110101",
						 "000001010100010001110010",
						 "000001010100010101101111",
						 "000001010100011001101100",
						 "000001010100011101101001",
						 "000001010100100001100110",
						 "000001010100100101100011",
						 "000001010100101001100000",
						 "000001010100101101011101",
						 "000001010100110001011010",
						 "000001010100110101010111",
						 "000001010100111001010100",
						 "000001010100111101010001",
						 "000001010110100100111100",
						 "000001010110101000111001",
						 "000001010110101100110110",
						 "000001010110110000110011",
						 "000001010110110100110000",
						 "000001010110111000101101",
						 "000001010110111100101010",
						 "000001010111000000100111",
						 "000001010111000100100100",
						 "000001010111001000100001",
						 "000001010111001100011110",
						 "000001010111010000011011",
						 "000001010111010100011000",
						 "000001010111011000010101",
						 "000001010111011100010010",
						 "000001010111100000001111",
						 "000001010110100100111100",
						 "000001010110101000111001",
						 "000001010110101100110110",
						 "000001010110110000110011",
						 "000001010110110100110000",
						 "000001010110111000101101",
						 "000001010110111100101010",
						 "000001010111000000100111",
						 "000001010111000100100100",
						 "000001010111001000100001",
						 "000001010111001100011110",
						 "000001010111010000011011",
						 "000001010111010100011000",
						 "000001010111011000010101",
						 "000001010111011100010010",
						 "000001010111100000001111",
						 "000001010110100100111100",
						 "000001010110101000111001",
						 "000001010110101100110110",
						 "000001010110110000110011",
						 "000001010110110100110000",
						 "000001010110111000101101",
						 "000001010110111100101010",
						 "000001010111000000100111",
						 "000001010111000100100100",
						 "000001010111001000100001",
						 "000001010111001100011110",
						 "000001010111010000011011",
						 "000001010111010100011000",
						 "000001010111011000010101",
						 "000001010111011100010010",
						 "000001010111100000001111",
						 "000001011001000111111010",
						 "000001011001001011110111",
						 "000001011001001111110100",
						 "000001011001010011110001",
						 "000001011001010111101110",
						 "000001011001011011101011",
						 "000001011001011111101000",
						 "000001011001100011100101",
						 "000001011001100111100010",
						 "000001011001101011011111",
						 "000001011001101111011100",
						 "000001011001110011011001",
						 "000001011001110111010110",
						 "000001011001111011010011",
						 "000001011001111111010000",
						 "000001011010000011001101",
						 "000001011001000111111010",
						 "000001011001001011110111",
						 "000001011001001111110100",
						 "000001011001010011110001",
						 "000001011001010111101110",
						 "000001011001011011101011",
						 "000001011001011111101000",
						 "000001011001100011100101",
						 "000001011001100111100010",
						 "000001011001101011011111",
						 "000001011001101111011100",
						 "000001011001110011011001",
						 "000001011001110111010110",
						 "000001011001111011010011",
						 "000001011001111111010000",
						 "000001011010000011001101",
						 "000001011001000111111010",
						 "000001011001001011110110",
						 "000001011001001111110010",
						 "000001011001010011101110",
						 "000001011001010111101010",
						 "000001011001011011100110",
						 "000001011001011111100010",
						 "000001011001100011011110",
						 "000001011001100111011010",
						 "000001011001101011010110",
						 "000001011001101111010010",
						 "000001011001110011001110",
						 "000001011001110111001010",
						 "000001011001111011000110",
						 "000001011001111111000010",
						 "000001011010000010111110",
						 "000001011011101010111000",
						 "000001011011101110110100",
						 "000001011011110010110000",
						 "000001011011110110101100",
						 "000001011011111010101000",
						 "000001011011111110100100",
						 "000001011100000010100000",
						 "000001011100000110011100",
						 "000001011100001010011000",
						 "000001011100001110010100",
						 "000001011100010010010000",
						 "000001011100010110001100",
						 "000001011100011010001000",
						 "000001011100011110000100",
						 "000001011100100010000000",
						 "000001011100100101111100",
						 "000001011011101010111000",
						 "000001011011101110110100",
						 "000001011011110010110000",
						 "000001011011110110101100",
						 "000001011011111010101000",
						 "000001011011111110100100",
						 "000001011100000010100000",
						 "000001011100000110011100",
						 "000001011100001010011000",
						 "000001011100001110010100",
						 "000001011100010010010000",
						 "000001011100010110001100",
						 "000001011100011010001000",
						 "000001011100011110000100",
						 "000001011100100010000000",
						 "000001011100100101111100",
						 "000001011110001101110110",
						 "000001011110010001110010",
						 "000001011110010101101110",
						 "000001011110011001101010",
						 "000001011110011101100110",
						 "000001011110100001100010",
						 "000001011110100101011110",
						 "000001011110101001011010",
						 "000001011110101101010110",
						 "000001011110110001010010",
						 "000001011110110101001110",
						 "000001011110111001001010",
						 "000001011110111101000110",
						 "000001011111000001000010",
						 "000001011111000100111110",
						 "000001011111001000111010",
						 "000001011110001101110110",
						 "000001011110010001110010",
						 "000001011110010101101110",
						 "000001011110011001101010",
						 "000001011110011101100110",
						 "000001011110100001100010",
						 "000001011110100101011110",
						 "000001011110101001011010",
						 "000001011110101101010110",
						 "000001011110110001010010",
						 "000001011110110101001110",
						 "000001011110111001001010",
						 "000001011110111101000110",
						 "000001011111000001000010",
						 "000001011111000100111110",
						 "000001011111001000111010",
						 "000001011110001101110110",
						 "000001011110010001110010",
						 "000001011110010101101110",
						 "000001011110011001101010",
						 "000001011110011101100110",
						 "000001011110100001100010",
						 "000001011110100101011110",
						 "000001011110101001011010",
						 "000001011110101101010110",
						 "000001011110110001010010",
						 "000001011110110101001110",
						 "000001011110111001001010",
						 "000001011110111101000110",
						 "000001011111000001000010",
						 "000001011111000100111110",
						 "000001011111001000111010",
						 "000001100000110000110100",
						 "000001100000110100110000",
						 "000001100000111000101100",
						 "000001100000111100101000",
						 "000001100001000000100100",
						 "000001100001000100100000",
						 "000001100001001000011100",
						 "000001100001001100011000",
						 "000001100001010000010100",
						 "000001100001010100010000",
						 "000001100001011000001100",
						 "000001100001011100001000",
						 "000001100001100000000100",
						 "000001100001100100000000",
						 "000001100001100111111100",
						 "000001100001101011111000",
						 "000001100000110000110100",
						 "000001100000110100110000",
						 "000001100000111000101100",
						 "000001100000111100101000",
						 "000001100001000000100100",
						 "000001100001000100100000",
						 "000001100001001000011100",
						 "000001100001001100011000",
						 "000001100001010000010100",
						 "000001100001010100010000",
						 "000001100001011000001100",
						 "000001100001011100001000",
						 "000001100001100000000100",
						 "000001100001100100000000",
						 "000001100001100111111100",
						 "000001100001101011111000",
						 "000001100011010011110010",
						 "000001100011010111101110",
						 "000001100011011011101010",
						 "000001100011011111100110",
						 "000001100011100011100010",
						 "000001100011100111011110",
						 "000001100011101011011010",
						 "000001100011101111010110",
						 "000001100011110011010010",
						 "000001100011110111001110",
						 "000001100011111011001010",
						 "000001100011111111000110",
						 "000001100100000011000010",
						 "000001100100000110111110",
						 "000001100100001010111010",
						 "000001100100001110110110",
						 "000001100011010011110010",
						 "000001100011010111101110",
						 "000001100011011011101010",
						 "000001100011011111100110",
						 "000001100011100011100010",
						 "000001100011100111011110",
						 "000001100011101011011010",
						 "000001100011101111010110",
						 "000001100011110011010010",
						 "000001100011110111001110",
						 "000001100011111011001010",
						 "000001100011111111000110",
						 "000001100100000011000010",
						 "000001100100000110111110",
						 "000001100100001010111010",
						 "000001100100001110110110",
						 "000001100011010011110010",
						 "000001100011010111101110",
						 "000001100011011011101010",
						 "000001100011011111100110",
						 "000001100011100011100010",
						 "000001100011100111011110",
						 "000001100011101011011010",
						 "000001100011101111010110",
						 "000001100011110011010010",
						 "000001100011110111001110",
						 "000001100011111011001010",
						 "000001100011111111000110",
						 "000001100100000011000010",
						 "000001100100000110111110",
						 "000001100100001010111010",
						 "000001100100001110110110",
						 "000001100101110110110000",
						 "000001100101111010101100",
						 "000001100101111110101000",
						 "000001100110000010100100",
						 "000001100110000110100000",
						 "000001100110001010011100",
						 "000001100110001110011000",
						 "000001100110010010010100",
						 "000001100110010110010000",
						 "000001100110011010001100",
						 "000001100110011110001000",
						 "000001100110100010000100",
						 "000001100110100110000000",
						 "000001100110101001111100",
						 "000001100110101101111000",
						 "000001100110110001110100",
						 "000001100101110110110000",
						 "000001100101111010101100",
						 "000001100101111110101000",
						 "000001100110000010100100",
						 "000001100110000110100000",
						 "000001100110001010011100",
						 "000001100110001110011000",
						 "000001100110010010010100",
						 "000001100110010110010000",
						 "000001100110011010001100",
						 "000001100110011110001000",
						 "000001100110100010000100",
						 "000001100110100110000000",
						 "000001100110101001111100",
						 "000001100110101101111000",
						 "000001100110110001110100",
						 "000001101000011001101110",
						 "000001101000011101101010",
						 "000001101000100001100110",
						 "000001101000100101100010",
						 "000001101000101001011110",
						 "000001101000101101011010",
						 "000001101000110001010110",
						 "000001101000110101010010",
						 "000001101000111001001110",
						 "000001101000111101001010",
						 "000001101001000001000110",
						 "000001101001000101000010",
						 "000001101001001000111110",
						 "000001101001001100111010",
						 "000001101001010000110110",
						 "000001101001010100110010",
						 "000001101000011001101110",
						 "000001101000011101101010",
						 "000001101000100001100110",
						 "000001101000100101100010",
						 "000001101000101001011110",
						 "000001101000101101011010",
						 "000001101000110001010110",
						 "000001101000110101010010",
						 "000001101000111001001110",
						 "000001101000111101001010",
						 "000001101001000001000110",
						 "000001101001000101000010",
						 "000001101001001000111110",
						 "000001101001001100111010",
						 "000001101001010000110110",
						 "000001101001010100110010",
						 "000001101000011001101110",
						 "000001101000011101101010",
						 "000001101000100001100110",
						 "000001101000100101100010",
						 "000001101000101001011110",
						 "000001101000101101011010",
						 "000001101000110001010110",
						 "000001101000110101010010",
						 "000001101000111001001110",
						 "000001101000111101001010",
						 "000001101001000001000110",
						 "000001101001000101000010",
						 "000001101001001000111110",
						 "000001101001001100111010",
						 "000001101001010000110110",
						 "000001101001010100110010",
						 "000001101010111100101100",
						 "000001101011000000101000",
						 "000001101011000100100100",
						 "000001101011001000100000",
						 "000001101011001100011100",
						 "000001101011010000011000",
						 "000001101011010100010100",
						 "000001101011011000010000",
						 "000001101011011100001100",
						 "000001101011100000001000",
						 "000001101011100100000100",
						 "000001101011101000000000",
						 "000001101011101011111100",
						 "000001101011101111111000",
						 "000001101011110011110100",
						 "000001101011110111110000",
						 "000001101010111100101100",
						 "000001101011000000100111",
						 "000001101011000100100010",
						 "000001101011001000011101",
						 "000001101011001100011000",
						 "000001101011010000010011",
						 "000001101011010100001110",
						 "000001101011011000001001",
						 "000001101011011100000100",
						 "000001101011011111111111",
						 "000001101011100011111010",
						 "000001101011100111110101",
						 "000001101011101011110000",
						 "000001101011101111101011",
						 "000001101011110011100110",
						 "000001101011110111100001",
						 "000001101010111100101100",
						 "000001101011000000100111",
						 "000001101011000100100010",
						 "000001101011001000011101",
						 "000001101011001100011000",
						 "000001101011010000010011",
						 "000001101011010100001110",
						 "000001101011011000001001",
						 "000001101011011100000100",
						 "000001101011011111111111",
						 "000001101011100011111010",
						 "000001101011100111110101",
						 "000001101011101011110000",
						 "000001101011101111101011",
						 "000001101011110011100110",
						 "000001101011110111100001",
						 "000001101101011111101010",
						 "000001101101100011100101",
						 "000001101101100111100000",
						 "000001101101101011011011",
						 "000001101101101111010110",
						 "000001101101110011010001",
						 "000001101101110111001100",
						 "000001101101111011000111",
						 "000001101101111111000010",
						 "000001101110000010111101",
						 "000001101110000110111000",
						 "000001101110001010110011",
						 "000001101110001110101110",
						 "000001101110010010101001",
						 "000001101110010110100100",
						 "000001101110011010011111",
						 "000001101101011111101010",
						 "000001101101100011100101",
						 "000001101101100111100000",
						 "000001101101101011011011",
						 "000001101101101111010110",
						 "000001101101110011010001",
						 "000001101101110111001100",
						 "000001101101111011000111",
						 "000001101101111111000010",
						 "000001101110000010111101",
						 "000001101110000110111000",
						 "000001101110001010110011",
						 "000001101110001110101110",
						 "000001101110010010101001",
						 "000001101110010110100100",
						 "000001101110011010011111",
						 "000001110000000010101000",
						 "000001110000000110100011",
						 "000001110000001010011110",
						 "000001110000001110011001",
						 "000001110000010010010100",
						 "000001110000010110001111",
						 "000001110000011010001010",
						 "000001110000011110000101",
						 "000001110000100010000000",
						 "000001110000100101111011",
						 "000001110000101001110110",
						 "000001110000101101110001",
						 "000001110000110001101100",
						 "000001110000110101100111",
						 "000001110000111001100010",
						 "000001110000111101011101",
						 "000001110000000010101000",
						 "000001110000000110100011",
						 "000001110000001010011110",
						 "000001110000001110011001",
						 "000001110000010010010100",
						 "000001110000010110001111",
						 "000001110000011010001010",
						 "000001110000011110000101",
						 "000001110000100010000000",
						 "000001110000100101111011",
						 "000001110000101001110110",
						 "000001110000101101110001",
						 "000001110000110001101100",
						 "000001110000110101100111",
						 "000001110000111001100010",
						 "000001110000111101011101",
						 "000001110000000010101000",
						 "000001110000000110100011",
						 "000001110000001010011110",
						 "000001110000001110011001",
						 "000001110000010010010100",
						 "000001110000010110001111",
						 "000001110000011010001010",
						 "000001110000011110000101",
						 "000001110000100010000000",
						 "000001110000100101111011",
						 "000001110000101001110110",
						 "000001110000101101110001",
						 "000001110000110001101100",
						 "000001110000110101100111",
						 "000001110000111001100010",
						 "000001110000111101011101",
						 "000001110010100101100110",
						 "000001110010101001100001",
						 "000001110010101101011100",
						 "000001110010110001010111",
						 "000001110010110101010010",
						 "000001110010111001001101",
						 "000001110010111101001000",
						 "000001110011000001000011",
						 "000001110011000100111110",
						 "000001110011001000111001",
						 "000001110011001100110100",
						 "000001110011010000101111",
						 "000001110011010100101010",
						 "000001110011011000100101",
						 "000001110011011100100000",
						 "000001110011100000011011",
						 "000001110010100101100110",
						 "000001110010101001100001",
						 "000001110010101101011100",
						 "000001110010110001010111",
						 "000001110010110101010010",
						 "000001110010111001001101",
						 "000001110010111101001000",
						 "000001110011000001000011",
						 "000001110011000100111110",
						 "000001110011001000111001",
						 "000001110011001100110100",
						 "000001110011010000101111",
						 "000001110011010100101010",
						 "000001110011011000100101",
						 "000001110011011100100000",
						 "000001110011100000011011",
						 "000001110101001000100100",
						 "000001110101001100011111",
						 "000001110101010000011010",
						 "000001110101010100010101",
						 "000001110101011000010000",
						 "000001110101011100001011",
						 "000001110101100000000110",
						 "000001110101100100000001",
						 "000001110101100111111100",
						 "000001110101101011110111",
						 "000001110101101111110010",
						 "000001110101110011101101",
						 "000001110101110111101000",
						 "000001110101111011100011",
						 "000001110101111111011110",
						 "000001110110000011011001",
						 "000001110101001000100100",
						 "000001110101001100011111",
						 "000001110101010000011010",
						 "000001110101010100010101",
						 "000001110101011000010000",
						 "000001110101011100001011",
						 "000001110101100000000110",
						 "000001110101100100000001",
						 "000001110101100111111100",
						 "000001110101101011110111",
						 "000001110101101111110010",
						 "000001110101110011101101",
						 "000001110101110111101000",
						 "000001110101111011100011",
						 "000001110101111111011110",
						 "000001110110000011011001",
						 "000001110101001000100100",
						 "000001110101001100011111",
						 "000001110101010000011010",
						 "000001110101010100010101",
						 "000001110101011000010000",
						 "000001110101011100001011",
						 "000001110101100000000110",
						 "000001110101100100000001",
						 "000001110101100111111100",
						 "000001110101101011110111",
						 "000001110101101111110010",
						 "000001110101110011101101",
						 "000001110101110111101000",
						 "000001110101111011100011",
						 "000001110101111111011110",
						 "000001110110000011011001",
						 "000001110111101011100010",
						 "000001110111101111011101",
						 "000001110111110011011000",
						 "000001110111110111010011",
						 "000001110111111011001110",
						 "000001110111111111001001",
						 "000001111000000011000100",
						 "000001111000000110111111",
						 "000001111000001010111010",
						 "000001111000001110110101",
						 "000001111000010010110000",
						 "000001111000010110101011",
						 "000001111000011010100110",
						 "000001111000011110100001",
						 "000001111000100010011100",
						 "000001111000100110010111",
						 "000001110111101011100010",
						 "000001110111101111011101",
						 "000001110111110011011000",
						 "000001110111110111010011",
						 "000001110111111011001110",
						 "000001110111111111001001",
						 "000001111000000011000100",
						 "000001111000000110111111",
						 "000001111000001010111010",
						 "000001111000001110110101",
						 "000001111000010010110000",
						 "000001111000010110101011",
						 "000001111000011010100110",
						 "000001111000011110100001",
						 "000001111000100010011100",
						 "000001111000100110010111",
						 "000001110111101011100010",
						 "000001110111101111011101",
						 "000001110111110011011000",
						 "000001110111110111010011",
						 "000001110111111011001110",
						 "000001110111111111001001",
						 "000001111000000011000100",
						 "000001111000000110111111",
						 "000001111000001010111010",
						 "000001111000001110110101",
						 "000001111000010010110000",
						 "000001111000010110101011",
						 "000001111000011010100110",
						 "000001111000011110100001",
						 "000001111000100010011100",
						 "000001111000100110010111",
						 "000001111010001110100000",
						 "000001111010010010011010",
						 "000001111010010110010100",
						 "000001111010011010001110",
						 "000001111010011110001000",
						 "000001111010100010000010",
						 "000001111010100101111100",
						 "000001111010101001110110",
						 "000001111010101101110000",
						 "000001111010110001101010",
						 "000001111010110101100100",
						 "000001111010111001011110",
						 "000001111010111101011000",
						 "000001111011000001010010",
						 "000001111011000101001100",
						 "000001111011001001000110",
						 "000001111010001110100000",
						 "000001111010010010011010",
						 "000001111010010110010100",
						 "000001111010011010001110",
						 "000001111010011110001000",
						 "000001111010100010000010",
						 "000001111010100101111100",
						 "000001111010101001110110",
						 "000001111010101101110000",
						 "000001111010110001101010",
						 "000001111010110101100100",
						 "000001111010111001011110",
						 "000001111010111101011000",
						 "000001111011000001010010",
						 "000001111011000101001100",
						 "000001111011001001000110",
						 "000001111100110001011110",
						 "000001111100110101011000",
						 "000001111100111001010010",
						 "000001111100111101001100",
						 "000001111101000001000110",
						 "000001111101000101000000",
						 "000001111101001000111010",
						 "000001111101001100110100",
						 "000001111101010000101110",
						 "000001111101010100101000",
						 "000001111101011000100010",
						 "000001111101011100011100",
						 "000001111101100000010110",
						 "000001111101100100010000",
						 "000001111101101000001010",
						 "000001111101101100000100",
						 "000001111100110001011110",
						 "000001111100110101011000",
						 "000001111100111001010010",
						 "000001111100111101001100",
						 "000001111101000001000110",
						 "000001111101000101000000",
						 "000001111101001000111010",
						 "000001111101001100110100",
						 "000001111101010000101110",
						 "000001111101010100101000",
						 "000001111101011000100010",
						 "000001111101011100011100",
						 "000001111101100000010110",
						 "000001111101100100010000",
						 "000001111101101000001010",
						 "000001111101101100000100",
						 "000001111100110001011110",
						 "000001111100110101011000",
						 "000001111100111001010010",
						 "000001111100111101001100",
						 "000001111101000001000110",
						 "000001111101000101000000",
						 "000001111101001000111010",
						 "000001111101001100110100",
						 "000001111101010000101110",
						 "000001111101010100101000",
						 "000001111101011000100010",
						 "000001111101011100011100",
						 "000001111101100000010110",
						 "000001111101100100010000",
						 "000001111101101000001010",
						 "000001111101101100000100",
						 "000001111111010100011100",
						 "000001111111011000010110",
						 "000001111111011100010000",
						 "000001111111100000001010",
						 "000001111111100100000100",
						 "000001111111100111111110",
						 "000001111111101011111000",
						 "000001111111101111110010",
						 "000001111111110011101100",
						 "000001111111110111100110",
						 "000001111111111011100000",
						 "000001111111111111011010",
						 "000010000000000011010100",
						 "000010000000000111001110",
						 "000010000000001011001000",
						 "000010000000001111000010",
						 "000001111111010100011100",
						 "000001111111011000010110",
						 "000001111111011100010000",
						 "000001111111100000001010",
						 "000001111111100100000100",
						 "000001111111100111111110",
						 "000001111111101011111000",
						 "000001111111101111110010",
						 "000001111111110011101100",
						 "000001111111110111100110",
						 "000001111111111011100000",
						 "000001111111111111011010",
						 "000010000000000011010100",
						 "000010000000000111001110",
						 "000010000000001011001000",
						 "000010000000001111000010",
						 "000010000001110111011010",
						 "000010000001111011010100",
						 "000010000001111111001110",
						 "000010000010000011001000",
						 "000010000010000111000010",
						 "000010000010001010111100",
						 "000010000010001110110110",
						 "000010000010010010110000",
						 "000010000010010110101010",
						 "000010000010011010100100",
						 "000010000010011110011110",
						 "000010000010100010011000",
						 "000010000010100110010010",
						 "000010000010101010001100",
						 "000010000010101110000110",
						 "000010000010110010000000",
						 "000010000001110111011010",
						 "000010000001111011010100",
						 "000010000001111111001110",
						 "000010000010000011001000",
						 "000010000010000111000010",
						 "000010000010001010111100",
						 "000010000010001110110110",
						 "000010000010010010110000",
						 "000010000010010110101010",
						 "000010000010011010100100",
						 "000010000010011110011110",
						 "000010000010100010011000",
						 "000010000010100110010010",
						 "000010000010101010001100",
						 "000010000010101110000110",
						 "000010000010110010000000",
						 "000010000001110111011010",
						 "000010000001111011010100",
						 "000010000001111111001110",
						 "000010000010000011001000",
						 "000010000010000111000010",
						 "000010000010001010111100",
						 "000010000010001110110110",
						 "000010000010010010110000",
						 "000010000010010110101010",
						 "000010000010011010100100",
						 "000010000010011110011110",
						 "000010000010100010011000",
						 "000010000010100110010010",
						 "000010000010101010001100",
						 "000010000010101110000110",
						 "000010000010110010000000",
						 "000010000100011010011000",
						 "000010000100011110010010",
						 "000010000100100010001100",
						 "000010000100100110000110",
						 "000010000100101010000000",
						 "000010000100101101111010",
						 "000010000100110001110100",
						 "000010000100110101101110",
						 "000010000100111001101000",
						 "000010000100111101100010",
						 "000010000101000001011100",
						 "000010000101000101010110",
						 "000010000101001001010000",
						 "000010000101001101001010",
						 "000010000101010001000100",
						 "000010000101010100111110",
						 "000010000100011010011000",
						 "000010000100011110010010",
						 "000010000100100010001100",
						 "000010000100100110000110",
						 "000010000100101010000000",
						 "000010000100101101111010",
						 "000010000100110001110100",
						 "000010000100110101101110",
						 "000010000100111001101000",
						 "000010000100111101100010",
						 "000010000101000001011100",
						 "000010000101000101010110",
						 "000010000101001001010000",
						 "000010000101001101001010",
						 "000010000101010001000100",
						 "000010000101010100111110",
						 "000010000100011010011000",
						 "000010000100011110010010",
						 "000010000100100010001100",
						 "000010000100100110000110",
						 "000010000100101010000000",
						 "000010000100101101111010",
						 "000010000100110001110100",
						 "000010000100110101101110",
						 "000010000100111001101000",
						 "000010000100111101100010",
						 "000010000101000001011100",
						 "000010000101000101010110",
						 "000010000101001001010000",
						 "000010000101001101001010",
						 "000010000101010001000100",
						 "000010000101010100111110",
						 "000010000110111101010110",
						 "000010000111000001001111",
						 "000010000111000101001000",
						 "000010000111001001000001",
						 "000010000111001100111010",
						 "000010000111010000110011",
						 "000010000111010100101100",
						 "000010000111011000100101",
						 "000010000111011100011110",
						 "000010000111100000010111",
						 "000010000111100100010000",
						 "000010000111101000001001",
						 "000010000111101100000010",
						 "000010000111101111111011",
						 "000010000111110011110100",
						 "000010000111110111101101",
						 "000010000110111101010110",
						 "000010000111000001001111",
						 "000010000111000101001000",
						 "000010000111001001000001",
						 "000010000111001100111010",
						 "000010000111010000110011",
						 "000010000111010100101100",
						 "000010000111011000100101",
						 "000010000111011100011110",
						 "000010000111100000010111",
						 "000010000111100100010000",
						 "000010000111101000001001",
						 "000010000111101100000010",
						 "000010000111101111111011",
						 "000010000111110011110100",
						 "000010000111110111101101",
						 "000010001001100000010100",
						 "000010001001100100001101",
						 "000010001001101000000110",
						 "000010001001101011111111",
						 "000010001001101111111000",
						 "000010001001110011110001",
						 "000010001001110111101010",
						 "000010001001111011100011",
						 "000010001001111111011100",
						 "000010001010000011010101",
						 "000010001010000111001110",
						 "000010001010001011000111",
						 "000010001010001111000000",
						 "000010001010010010111001",
						 "000010001010010110110010",
						 "000010001010011010101011",
						 "000010001001100000010100",
						 "000010001001100100001101",
						 "000010001001101000000110",
						 "000010001001101011111111",
						 "000010001001101111111000",
						 "000010001001110011110001",
						 "000010001001110111101010",
						 "000010001001111011100011",
						 "000010001001111111011100",
						 "000010001010000011010101",
						 "000010001010000111001110",
						 "000010001010001011000111",
						 "000010001010001111000000",
						 "000010001010010010111001",
						 "000010001010010110110010",
						 "000010001010011010101011",
						 "000010001001100000010100",
						 "000010001001100100001101",
						 "000010001001101000000110",
						 "000010001001101011111111",
						 "000010001001101111111000",
						 "000010001001110011110001",
						 "000010001001110111101010",
						 "000010001001111011100011",
						 "000010001001111111011100",
						 "000010001010000011010101",
						 "000010001010000111001110",
						 "000010001010001011000111",
						 "000010001010001111000000",
						 "000010001010010010111001",
						 "000010001010010110110010",
						 "000010001010011010101011",
						 "000010001100000011010010",
						 "000010001100000111001011",
						 "000010001100001011000100",
						 "000010001100001110111101",
						 "000010001100010010110110",
						 "000010001100010110101111",
						 "000010001100011010101000",
						 "000010001100011110100001",
						 "000010001100100010011010",
						 "000010001100100110010011",
						 "000010001100101010001100",
						 "000010001100101110000101",
						 "000010001100110001111110",
						 "000010001100110101110111",
						 "000010001100111001110000",
						 "000010001100111101101001",
						 "000010001100000011010010",
						 "000010001100000111001011",
						 "000010001100001011000100",
						 "000010001100001110111101",
						 "000010001100010010110110",
						 "000010001100010110101111",
						 "000010001100011010101000",
						 "000010001100011110100001",
						 "000010001100100010011010",
						 "000010001100100110010011",
						 "000010001100101010001100",
						 "000010001100101110000101",
						 "000010001100110001111110",
						 "000010001100110101110111",
						 "000010001100111001110000",
						 "000010001100111101101001",
						 "000010001100000011010010",
						 "000010001100000111001011",
						 "000010001100001011000100",
						 "000010001100001110111101",
						 "000010001100010010110110",
						 "000010001100010110101111",
						 "000010001100011010101000",
						 "000010001100011110100001",
						 "000010001100100010011010",
						 "000010001100100110010011",
						 "000010001100101010001100",
						 "000010001100101110000101",
						 "000010001100110001111110",
						 "000010001100110101110111",
						 "000010001100111001110000",
						 "000010001100111101101001",
						 "000010001110100110010000",
						 "000010001110101010001001",
						 "000010001110101110000010",
						 "000010001110110001111011",
						 "000010001110110101110100",
						 "000010001110111001101101",
						 "000010001110111101100110",
						 "000010001111000001011111",
						 "000010001111000101011000",
						 "000010001111001001010001",
						 "000010001111001101001010",
						 "000010001111010001000011",
						 "000010001111010100111100",
						 "000010001111011000110101",
						 "000010001111011100101110",
						 "000010001111100000100111",
						 "000010001110100110010000",
						 "000010001110101010001001",
						 "000010001110101110000010",
						 "000010001110110001111011",
						 "000010001110110101110100",
						 "000010001110111001101101",
						 "000010001110111101100110",
						 "000010001111000001011111",
						 "000010001111000101011000",
						 "000010001111001001010001",
						 "000010001111001101001010",
						 "000010001111010001000011",
						 "000010001111010100111100",
						 "000010001111011000110101",
						 "000010001111011100101110",
						 "000010001111100000100111",
						 "000010010001001001001110",
						 "000010010001001101000111",
						 "000010010001010001000000",
						 "000010010001010100111001",
						 "000010010001011000110010",
						 "000010010001011100101011",
						 "000010010001100000100100",
						 "000010010001100100011101",
						 "000010010001101000010110",
						 "000010010001101100001111",
						 "000010010001110000001000",
						 "000010010001110100000001",
						 "000010010001110111111010",
						 "000010010001111011110011",
						 "000010010001111111101100",
						 "000010010010000011100101",
						 "000010010001001001001110",
						 "000010010001001101000111",
						 "000010010001010001000000",
						 "000010010001010100111001",
						 "000010010001011000110010",
						 "000010010001011100101011",
						 "000010010001100000100100",
						 "000010010001100100011101",
						 "000010010001101000010110",
						 "000010010001101100001111",
						 "000010010001110000001000",
						 "000010010001110100000001",
						 "000010010001110111111010",
						 "000010010001111011110011",
						 "000010010001111111101100",
						 "000010010010000011100101",
						 "000010010001001001001110",
						 "000010010001001101000110",
						 "000010010001010000111110",
						 "000010010001010100110110",
						 "000010010001011000101110",
						 "000010010001011100100110",
						 "000010010001100000011110",
						 "000010010001100100010110",
						 "000010010001101000001110",
						 "000010010001101100000110",
						 "000010010001101111111110",
						 "000010010001110011110110",
						 "000010010001110111101110",
						 "000010010001111011100110",
						 "000010010001111111011110",
						 "000010010010000011010110",
						 "000010010011101100001100",
						 "000010010011110000000100",
						 "000010010011110011111100",
						 "000010010011110111110100",
						 "000010010011111011101100",
						 "000010010011111111100100",
						 "000010010100000011011100",
						 "000010010100000111010100",
						 "000010010100001011001100",
						 "000010010100001111000100",
						 "000010010100010010111100",
						 "000010010100010110110100",
						 "000010010100011010101100",
						 "000010010100011110100100",
						 "000010010100100010011100",
						 "000010010100100110010100",
						 "000010010011101100001100",
						 "000010010011110000000100",
						 "000010010011110011111100",
						 "000010010011110111110100",
						 "000010010011111011101100",
						 "000010010011111111100100",
						 "000010010100000011011100",
						 "000010010100000111010100",
						 "000010010100001011001100",
						 "000010010100001111000100",
						 "000010010100010010111100",
						 "000010010100010110110100",
						 "000010010100011010101100",
						 "000010010100011110100100",
						 "000010010100100010011100",
						 "000010010100100110010100",
						 "000010010110001111001010",
						 "000010010110010011000010",
						 "000010010110010110111010",
						 "000010010110011010110010",
						 "000010010110011110101010",
						 "000010010110100010100010",
						 "000010010110100110011010",
						 "000010010110101010010010",
						 "000010010110101110001010",
						 "000010010110110010000010",
						 "000010010110110101111010",
						 "000010010110111001110010",
						 "000010010110111101101010",
						 "000010010111000001100010",
						 "000010010111000101011010",
						 "000010010111001001010010",
						 "000010010110001111001010",
						 "000010010110010011000010",
						 "000010010110010110111010",
						 "000010010110011010110010",
						 "000010010110011110101010",
						 "000010010110100010100010",
						 "000010010110100110011010",
						 "000010010110101010010010",
						 "000010010110101110001010",
						 "000010010110110010000010",
						 "000010010110110101111010",
						 "000010010110111001110010",
						 "000010010110111101101010",
						 "000010010111000001100010",
						 "000010010111000101011010",
						 "000010010111001001010010",
						 "000010010110001111001010",
						 "000010010110010011000010",
						 "000010010110010110111010",
						 "000010010110011010110010",
						 "000010010110011110101010",
						 "000010010110100010100010",
						 "000010010110100110011010",
						 "000010010110101010010010",
						 "000010010110101110001010",
						 "000010010110110010000010",
						 "000010010110110101111010",
						 "000010010110111001110010",
						 "000010010110111101101010",
						 "000010010111000001100010",
						 "000010010111000101011010",
						 "000010010111001001010010",
						 "000010011000110010001000",
						 "000010011000110110000000",
						 "000010011000111001111000",
						 "000010011000111101110000",
						 "000010011001000001101000",
						 "000010011001000101100000",
						 "000010011001001001011000",
						 "000010011001001101010000",
						 "000010011001010001001000",
						 "000010011001010101000000",
						 "000010011001011000111000",
						 "000010011001011100110000",
						 "000010011001100000101000",
						 "000010011001100100100000",
						 "000010011001101000011000",
						 "000010011001101100010000",
						 "000010011000110010001000",
						 "000010011000110110000000",
						 "000010011000111001111000",
						 "000010011000111101110000",
						 "000010011001000001101000",
						 "000010011001000101100000",
						 "000010011001001001011000",
						 "000010011001001101010000",
						 "000010011001010001001000",
						 "000010011001010101000000",
						 "000010011001011000111000",
						 "000010011001011100110000",
						 "000010011001100000101000",
						 "000010011001100100100000",
						 "000010011001101000011000",
						 "000010011001101100010000",
						 "000010011000110010001000",
						 "000010011000110110000000",
						 "000010011000111001111000",
						 "000010011000111101110000",
						 "000010011001000001101000",
						 "000010011001000101100000",
						 "000010011001001001011000",
						 "000010011001001101010000",
						 "000010011001010001001000",
						 "000010011001010101000000",
						 "000010011001011000111000",
						 "000010011001011100110000",
						 "000010011001100000101000",
						 "000010011001100100100000",
						 "000010011001101000011000",
						 "000010011001101100010000",
						 "000010011011010101000110",
						 "000010011011011000111110",
						 "000010011011011100110110",
						 "000010011011100000101110",
						 "000010011011100100100110",
						 "000010011011101000011110",
						 "000010011011101100010110",
						 "000010011011110000001110",
						 "000010011011110100000110",
						 "000010011011110111111110",
						 "000010011011111011110110",
						 "000010011011111111101110",
						 "000010011100000011100110",
						 "000010011100000111011110",
						 "000010011100001011010110",
						 "000010011100001111001110",
						 "000010011011010101000110",
						 "000010011011011000111101",
						 "000010011011011100110100",
						 "000010011011100000101011",
						 "000010011011100100100010",
						 "000010011011101000011001",
						 "000010011011101100010000",
						 "000010011011110000000111",
						 "000010011011110011111110",
						 "000010011011110111110101",
						 "000010011011111011101100",
						 "000010011011111111100011",
						 "000010011100000011011010",
						 "000010011100000111010001",
						 "000010011100001011001000",
						 "000010011100001110111111",
						 "000010011101111000000100",
						 "000010011101111011111011",
						 "000010011101111111110010",
						 "000010011110000011101001",
						 "000010011110000111100000",
						 "000010011110001011010111",
						 "000010011110001111001110",
						 "000010011110010011000101",
						 "000010011110010110111100",
						 "000010011110011010110011",
						 "000010011110011110101010",
						 "000010011110100010100001",
						 "000010011110100110011000",
						 "000010011110101010001111",
						 "000010011110101110000110",
						 "000010011110110001111101",
						 "000010011101111000000100",
						 "000010011101111011111011",
						 "000010011101111111110010",
						 "000010011110000011101001",
						 "000010011110000111100000",
						 "000010011110001011010111",
						 "000010011110001111001110",
						 "000010011110010011000101",
						 "000010011110010110111100",
						 "000010011110011010110011",
						 "000010011110011110101010",
						 "000010011110100010100001",
						 "000010011110100110011000",
						 "000010011110101010001111",
						 "000010011110101110000110",
						 "000010011110110001111101",
						 "000010011101111000000100",
						 "000010011101111011111011",
						 "000010011101111111110010",
						 "000010011110000011101001",
						 "000010011110000111100000",
						 "000010011110001011010111",
						 "000010011110001111001110",
						 "000010011110010011000101",
						 "000010011110010110111100",
						 "000010011110011010110011",
						 "000010011110011110101010",
						 "000010011110100010100001",
						 "000010011110100110011000",
						 "000010011110101010001111",
						 "000010011110101110000110",
						 "000010011110110001111101",
						 "000010100000011011000010",
						 "000010100000011110111001",
						 "000010100000100010110000",
						 "000010100000100110100111",
						 "000010100000101010011110",
						 "000010100000101110010101",
						 "000010100000110010001100",
						 "000010100000110110000011",
						 "000010100000111001111010",
						 "000010100000111101110001",
						 "000010100001000001101000",
						 "000010100001000101011111",
						 "000010100001001001010110",
						 "000010100001001101001101",
						 "000010100001010001000100",
						 "000010100001010100111011",
						 "000010100000011011000010",
						 "000010100000011110111001",
						 "000010100000100010110000",
						 "000010100000100110100111",
						 "000010100000101010011110",
						 "000010100000101110010101",
						 "000010100000110010001100",
						 "000010100000110110000011",
						 "000010100000111001111010",
						 "000010100000111101110001",
						 "000010100001000001101000",
						 "000010100001000101011111",
						 "000010100001001001010110",
						 "000010100001001101001101",
						 "000010100001010001000100",
						 "000010100001010100111011",
						 "000010100000011011000010",
						 "000010100000011110111001",
						 "000010100000100010110000",
						 "000010100000100110100111",
						 "000010100000101010011110",
						 "000010100000101110010101",
						 "000010100000110010001100",
						 "000010100000110110000011",
						 "000010100000111001111010",
						 "000010100000111101110001",
						 "000010100001000001101000",
						 "000010100001000101011111",
						 "000010100001001001010110",
						 "000010100001001101001101",
						 "000010100001010001000100",
						 "000010100001010100111011",
						 "000010100010111110000000",
						 "000010100011000001110111",
						 "000010100011000101101110",
						 "000010100011001001100101",
						 "000010100011001101011100",
						 "000010100011010001010011",
						 "000010100011010101001010",
						 "000010100011011001000001",
						 "000010100011011100111000",
						 "000010100011100000101111",
						 "000010100011100100100110",
						 "000010100011101000011101",
						 "000010100011101100010100",
						 "000010100011110000001011",
						 "000010100011110100000010",
						 "000010100011110111111001",
						 "000010100010111110000000",
						 "000010100011000001110111",
						 "000010100011000101101110",
						 "000010100011001001100101",
						 "000010100011001101011100",
						 "000010100011010001010011",
						 "000010100011010101001010",
						 "000010100011011001000001",
						 "000010100011011100111000",
						 "000010100011100000101111",
						 "000010100011100100100110",
						 "000010100011101000011101",
						 "000010100011101100010100",
						 "000010100011110000001011",
						 "000010100011110100000010",
						 "000010100011110111111001",
						 "000010100101100000111110",
						 "000010100101100100110101",
						 "000010100101101000101100",
						 "000010100101101100100011",
						 "000010100101110000011010",
						 "000010100101110100010001",
						 "000010100101111000001000",
						 "000010100101111011111111",
						 "000010100101111111110110",
						 "000010100110000011101101",
						 "000010100110000111100100",
						 "000010100110001011011011",
						 "000010100110001111010010",
						 "000010100110010011001001",
						 "000010100110010111000000",
						 "000010100110011010110111",
						 "000010100101100000111110",
						 "000010100101100100110101",
						 "000010100101101000101100",
						 "000010100101101100100011",
						 "000010100101110000011010",
						 "000010100101110100010001",
						 "000010100101111000001000",
						 "000010100101111011111111",
						 "000010100101111111110110",
						 "000010100110000011101101",
						 "000010100110000111100100",
						 "000010100110001011011011",
						 "000010100110001111010010",
						 "000010100110010011001001",
						 "000010100110010111000000",
						 "000010100110011010110111",
						 "000010100101100000111110",
						 "000010100101100100110100",
						 "000010100101101000101010",
						 "000010100101101100100000",
						 "000010100101110000010110",
						 "000010100101110100001100",
						 "000010100101111000000010",
						 "000010100101111011111000",
						 "000010100101111111101110",
						 "000010100110000011100100",
						 "000010100110000111011010",
						 "000010100110001011010000",
						 "000010100110001111000110",
						 "000010100110010010111100",
						 "000010100110010110110010",
						 "000010100110011010101000",
						 "000010101000000011111100",
						 "000010101000000111110010",
						 "000010101000001011101000",
						 "000010101000001111011110",
						 "000010101000010011010100",
						 "000010101000010111001010",
						 "000010101000011011000000",
						 "000010101000011110110110",
						 "000010101000100010101100",
						 "000010101000100110100010",
						 "000010101000101010011000",
						 "000010101000101110001110",
						 "000010101000110010000100",
						 "000010101000110101111010",
						 "000010101000111001110000",
						 "000010101000111101100110",
						 "000010101000000011111100",
						 "000010101000000111110010",
						 "000010101000001011101000",
						 "000010101000001111011110",
						 "000010101000010011010100",
						 "000010101000010111001010",
						 "000010101000011011000000",
						 "000010101000011110110110",
						 "000010101000100010101100",
						 "000010101000100110100010",
						 "000010101000101010011000",
						 "000010101000101110001110",
						 "000010101000110010000100",
						 "000010101000110101111010",
						 "000010101000111001110000",
						 "000010101000111101100110",
						 "000010101010100110111010",
						 "000010101010101010110000",
						 "000010101010101110100110",
						 "000010101010110010011100",
						 "000010101010110110010010",
						 "000010101010111010001000",
						 "000010101010111101111110",
						 "000010101011000001110100",
						 "000010101011000101101010",
						 "000010101011001001100000",
						 "000010101011001101010110",
						 "000010101011010001001100",
						 "000010101011010101000010",
						 "000010101011011000111000",
						 "000010101011011100101110",
						 "000010101011100000100100",
						 "000010101010100110111010",
						 "000010101010101010110000",
						 "000010101010101110100110",
						 "000010101010110010011100",
						 "000010101010110110010010",
						 "000010101010111010001000",
						 "000010101010111101111110",
						 "000010101011000001110100",
						 "000010101011000101101010",
						 "000010101011001001100000",
						 "000010101011001101010110",
						 "000010101011010001001100",
						 "000010101011010101000010",
						 "000010101011011000111000",
						 "000010101011011100101110",
						 "000010101011100000100100",
						 "000010101010100110111010",
						 "000010101010101010110000",
						 "000010101010101110100110",
						 "000010101010110010011100",
						 "000010101010110110010010",
						 "000010101010111010001000",
						 "000010101010111101111110",
						 "000010101011000001110100",
						 "000010101011000101101010",
						 "000010101011001001100000",
						 "000010101011001101010110",
						 "000010101011010001001100",
						 "000010101011010101000010",
						 "000010101011011000111000",
						 "000010101011011100101110",
						 "000010101011100000100100",
						 "000010101101001001111000",
						 "000010101101001101101110",
						 "000010101101010001100100",
						 "000010101101010101011010",
						 "000010101101011001010000",
						 "000010101101011101000110",
						 "000010101101100000111100",
						 "000010101101100100110010",
						 "000010101101101000101000",
						 "000010101101101100011110",
						 "000010101101110000010100",
						 "000010101101110100001010",
						 "000010101101111000000000",
						 "000010101101111011110110",
						 "000010101101111111101100",
						 "000010101110000011100010",
						 "000010101101001001111000",
						 "000010101101001101101110",
						 "000010101101010001100100",
						 "000010101101010101011010",
						 "000010101101011001010000",
						 "000010101101011101000110",
						 "000010101101100000111100",
						 "000010101101100100110010",
						 "000010101101101000101000",
						 "000010101101101100011110",
						 "000010101101110000010100",
						 "000010101101110100001010",
						 "000010101101111000000000",
						 "000010101101111011110110",
						 "000010101101111111101100",
						 "000010101110000011100010",
						 "000010101101001001111000",
						 "000010101101001101101110",
						 "000010101101010001100100",
						 "000010101101010101011010",
						 "000010101101011001010000",
						 "000010101101011101000110",
						 "000010101101100000111100",
						 "000010101101100100110010",
						 "000010101101101000101000",
						 "000010101101101100011110",
						 "000010101101110000010100",
						 "000010101101110100001010",
						 "000010101101111000000000",
						 "000010101101111011110110",
						 "000010101101111111101100",
						 "000010101110000011100010",
						 "000010101111101100110110",
						 "000010101111110000101011",
						 "000010101111110100100000",
						 "000010101111111000010101",
						 "000010101111111100001010",
						 "000010101111111111111111",
						 "000010110000000011110100",
						 "000010110000000111101001",
						 "000010110000001011011110",
						 "000010110000001111010011",
						 "000010110000010011001000",
						 "000010110000010110111101",
						 "000010110000011010110010",
						 "000010110000011110100111",
						 "000010110000100010011100",
						 "000010110000100110010001",
						 "000010101111101100110110",
						 "000010101111110000101011",
						 "000010101111110100100000",
						 "000010101111111000010101",
						 "000010101111111100001010",
						 "000010101111111111111111",
						 "000010110000000011110100",
						 "000010110000000111101001",
						 "000010110000001011011110",
						 "000010110000001111010011",
						 "000010110000010011001000",
						 "000010110000010110111101",
						 "000010110000011010110010",
						 "000010110000011110100111",
						 "000010110000100010011100",
						 "000010110000100110010001",
						 "000010110010001111110100",
						 "000010110010010011101001",
						 "000010110010010111011110",
						 "000010110010011011010011",
						 "000010110010011111001000",
						 "000010110010100010111101",
						 "000010110010100110110010",
						 "000010110010101010100111",
						 "000010110010101110011100",
						 "000010110010110010010001",
						 "000010110010110110000110",
						 "000010110010111001111011",
						 "000010110010111101110000",
						 "000010110011000001100101",
						 "000010110011000101011010",
						 "000010110011001001001111",
						 "000010110010001111110100",
						 "000010110010010011101001",
						 "000010110010010111011110",
						 "000010110010011011010011",
						 "000010110010011111001000",
						 "000010110010100010111101",
						 "000010110010100110110010",
						 "000010110010101010100111",
						 "000010110010101110011100",
						 "000010110010110010010001",
						 "000010110010110110000110",
						 "000010110010111001111011",
						 "000010110010111101110000",
						 "000010110011000001100101",
						 "000010110011000101011010",
						 "000010110011001001001111",
						 "000010110010001111110100",
						 "000010110010010011101001",
						 "000010110010010111011110",
						 "000010110010011011010011",
						 "000010110010011111001000",
						 "000010110010100010111101",
						 "000010110010100110110010",
						 "000010110010101010100111",
						 "000010110010101110011100",
						 "000010110010110010010001",
						 "000010110010110110000110",
						 "000010110010111001111011",
						 "000010110010111101110000",
						 "000010110011000001100101",
						 "000010110011000101011010",
						 "000010110011001001001111",
						 "000010110100110010110010",
						 "000010110100110110100111",
						 "000010110100111010011100",
						 "000010110100111110010001",
						 "000010110101000010000110",
						 "000010110101000101111011",
						 "000010110101001001110000",
						 "000010110101001101100101",
						 "000010110101010001011010",
						 "000010110101010101001111",
						 "000010110101011001000100",
						 "000010110101011100111001",
						 "000010110101100000101110",
						 "000010110101100100100011",
						 "000010110101101000011000",
						 "000010110101101100001101",
						 "000010110100110010110010",
						 "000010110100110110100111",
						 "000010110100111010011100",
						 "000010110100111110010001",
						 "000010110101000010000110",
						 "000010110101000101111011",
						 "000010110101001001110000",
						 "000010110101001101100101",
						 "000010110101010001011010",
						 "000010110101010101001111",
						 "000010110101011001000100",
						 "000010110101011100111001",
						 "000010110101100000101110",
						 "000010110101100100100011",
						 "000010110101101000011000",
						 "000010110101101100001101",
						 "000010110100110010110010",
						 "000010110100110110100111",
						 "000010110100111010011100",
						 "000010110100111110010001",
						 "000010110101000010000110",
						 "000010110101000101111011",
						 "000010110101001001110000",
						 "000010110101001101100101",
						 "000010110101010001011010",
						 "000010110101010101001111",
						 "000010110101011001000100",
						 "000010110101011100111001",
						 "000010110101100000101110",
						 "000010110101100100100011",
						 "000010110101101000011000",
						 "000010110101101100001101",
						 "000010110111010101110000",
						 "000010110111011001100101",
						 "000010110111011101011010",
						 "000010110111100001001111",
						 "000010110111100101000100",
						 "000010110111101000111001",
						 "000010110111101100101110",
						 "000010110111110000100011",
						 "000010110111110100011000",
						 "000010110111111000001101",
						 "000010110111111100000010",
						 "000010110111111111110111",
						 "000010111000000011101100",
						 "000010111000000111100001",
						 "000010111000001011010110",
						 "000010111000001111001011",
						 "000010110111010101110000",
						 "000010110111011001100101",
						 "000010110111011101011010",
						 "000010110111100001001111",
						 "000010110111100101000100",
						 "000010110111101000111001",
						 "000010110111101100101110",
						 "000010110111110000100011",
						 "000010110111110100011000",
						 "000010110111111000001101",
						 "000010110111111100000010",
						 "000010110111111111110111",
						 "000010111000000011101100",
						 "000010111000000111100001",
						 "000010111000001011010110",
						 "000010111000001111001011",
						 "000010111001111000101110",
						 "000010111001111100100010",
						 "000010111010000000010110",
						 "000010111010000100001010",
						 "000010111010000111111110",
						 "000010111010001011110010",
						 "000010111010001111100110",
						 "000010111010010011011010",
						 "000010111010010111001110",
						 "000010111010011011000010",
						 "000010111010011110110110",
						 "000010111010100010101010",
						 "000010111010100110011110",
						 "000010111010101010010010",
						 "000010111010101110000110",
						 "000010111010110001111010",
						 "000010111001111000101110",
						 "000010111001111100100010",
						 "000010111010000000010110",
						 "000010111010000100001010",
						 "000010111010000111111110",
						 "000010111010001011110010",
						 "000010111010001111100110",
						 "000010111010010011011010",
						 "000010111010010111001110",
						 "000010111010011011000010",
						 "000010111010011110110110",
						 "000010111010100010101010",
						 "000010111010100110011110",
						 "000010111010101010010010",
						 "000010111010101110000110",
						 "000010111010110001111010",
						 "000010111001111000101110",
						 "000010111001111100100010",
						 "000010111010000000010110",
						 "000010111010000100001010",
						 "000010111010000111111110",
						 "000010111010001011110010",
						 "000010111010001111100110",
						 "000010111010010011011010",
						 "000010111010010111001110",
						 "000010111010011011000010",
						 "000010111010011110110110",
						 "000010111010100010101010",
						 "000010111010100110011110",
						 "000010111010101010010010",
						 "000010111010101110000110",
						 "000010111010110001111010",
						 "000010111100011011101100",
						 "000010111100011111100000",
						 "000010111100100011010100",
						 "000010111100100111001000",
						 "000010111100101010111100",
						 "000010111100101110110000",
						 "000010111100110010100100",
						 "000010111100110110011000",
						 "000010111100111010001100",
						 "000010111100111110000000",
						 "000010111101000001110100",
						 "000010111101000101101000",
						 "000010111101001001011100",
						 "000010111101001101010000",
						 "000010111101010001000100",
						 "000010111101010100111000",
						 "000010111100011011101100",
						 "000010111100011111100000",
						 "000010111100100011010100",
						 "000010111100100111001000",
						 "000010111100101010111100",
						 "000010111100101110110000",
						 "000010111100110010100100",
						 "000010111100110110011000",
						 "000010111100111010001100",
						 "000010111100111110000000",
						 "000010111101000001110100",
						 "000010111101000101101000",
						 "000010111101001001011100",
						 "000010111101001101010000",
						 "000010111101010001000100",
						 "000010111101010100111000",
						 "000010111100011011101100",
						 "000010111100011111100000",
						 "000010111100100011010100",
						 "000010111100100111001000",
						 "000010111100101010111100",
						 "000010111100101110110000",
						 "000010111100110010100100",
						 "000010111100110110011000",
						 "000010111100111010001100",
						 "000010111100111110000000",
						 "000010111101000001110100",
						 "000010111101000101101000",
						 "000010111101001001011100",
						 "000010111101001101010000",
						 "000010111101010001000100",
						 "000010111101010100111000",
						 "000010111110111110101010",
						 "000010111111000010011110",
						 "000010111111000110010010",
						 "000010111111001010000110",
						 "000010111111001101111010",
						 "000010111111010001101110",
						 "000010111111010101100010",
						 "000010111111011001010110",
						 "000010111111011101001010",
						 "000010111111100000111110",
						 "000010111111100100110010",
						 "000010111111101000100110",
						 "000010111111101100011010",
						 "000010111111110000001110",
						 "000010111111110100000010",
						 "000010111111110111110110",
						 "000010111110111110101010",
						 "000010111111000010011110",
						 "000010111111000110010010",
						 "000010111111001010000110",
						 "000010111111001101111010",
						 "000010111111010001101110",
						 "000010111111010101100010",
						 "000010111111011001010110",
						 "000010111111011101001010",
						 "000010111111100000111110",
						 "000010111111100100110010",
						 "000010111111101000100110",
						 "000010111111101100011010",
						 "000010111111110000001110",
						 "000010111111110100000010",
						 "000010111111110111110110",
						 "000011000001100001101000",
						 "000011000001100101011100",
						 "000011000001101001010000",
						 "000011000001101101000100",
						 "000011000001110000111000",
						 "000011000001110100101100",
						 "000011000001111000100000",
						 "000011000001111100010100",
						 "000011000010000000001000",
						 "000011000010000011111100",
						 "000011000010000111110000",
						 "000011000010001011100100",
						 "000011000010001111011000",
						 "000011000010010011001100",
						 "000011000010010111000000",
						 "000011000010011010110100",
						 "000011000001100001101000",
						 "000011000001100101011011",
						 "000011000001101001001110",
						 "000011000001101101000001",
						 "000011000001110000110100",
						 "000011000001110100100111",
						 "000011000001111000011010",
						 "000011000001111100001101",
						 "000011000010000000000000",
						 "000011000010000011110011",
						 "000011000010000111100110",
						 "000011000010001011011001",
						 "000011000010001111001100",
						 "000011000010010010111111",
						 "000011000010010110110010",
						 "000011000010011010100101",
						 "000011000001100001101000",
						 "000011000001100101011011",
						 "000011000001101001001110",
						 "000011000001101101000001",
						 "000011000001110000110100",
						 "000011000001110100100111",
						 "000011000001111000011010",
						 "000011000001111100001101",
						 "000011000010000000000000",
						 "000011000010000011110011",
						 "000011000010000111100110",
						 "000011000010001011011001",
						 "000011000010001111001100",
						 "000011000010010010111111",
						 "000011000010010110110010",
						 "000011000010011010100101",
						 "000011000100000100100110",
						 "000011000100001000011001",
						 "000011000100001100001100",
						 "000011000100001111111111",
						 "000011000100010011110010",
						 "000011000100010111100101",
						 "000011000100011011011000",
						 "000011000100011111001011",
						 "000011000100100010111110",
						 "000011000100100110110001",
						 "000011000100101010100100",
						 "000011000100101110010111",
						 "000011000100110010001010",
						 "000011000100110101111101",
						 "000011000100111001110000",
						 "000011000100111101100011",
						 "000011000100000100100110",
						 "000011000100001000011001",
						 "000011000100001100001100",
						 "000011000100001111111111",
						 "000011000100010011110010",
						 "000011000100010111100101",
						 "000011000100011011011000",
						 "000011000100011111001011",
						 "000011000100100010111110",
						 "000011000100100110110001",
						 "000011000100101010100100",
						 "000011000100101110010111",
						 "000011000100110010001010",
						 "000011000100110101111101",
						 "000011000100111001110000",
						 "000011000100111101100011",
						 "000011000100000100100110",
						 "000011000100001000011001",
						 "000011000100001100001100",
						 "000011000100001111111111",
						 "000011000100010011110010",
						 "000011000100010111100101",
						 "000011000100011011011000",
						 "000011000100011111001011",
						 "000011000100100010111110",
						 "000011000100100110110001",
						 "000011000100101010100100",
						 "000011000100101110010111",
						 "000011000100110010001010",
						 "000011000100110101111101",
						 "000011000100111001110000",
						 "000011000100111101100011",
						 "000011000110100111100100",
						 "000011000110101011010111",
						 "000011000110101111001010",
						 "000011000110110010111101",
						 "000011000110110110110000",
						 "000011000110111010100011",
						 "000011000110111110010110",
						 "000011000111000010001001",
						 "000011000111000101111100",
						 "000011000111001001101111",
						 "000011000111001101100010",
						 "000011000111010001010101",
						 "000011000111010101001000",
						 "000011000111011000111011",
						 "000011000111011100101110",
						 "000011000111100000100001",
						 "000011000110100111100100",
						 "000011000110101011010111",
						 "000011000110101111001010",
						 "000011000110110010111101",
						 "000011000110110110110000",
						 "000011000110111010100011",
						 "000011000110111110010110",
						 "000011000111000010001001",
						 "000011000111000101111100",
						 "000011000111001001101111",
						 "000011000111001101100010",
						 "000011000111010001010101",
						 "000011000111010101001000",
						 "000011000111011000111011",
						 "000011000111011100101110",
						 "000011000111100000100001",
						 "000011001001001010100010",
						 "000011001001001110010101",
						 "000011001001010010001000",
						 "000011001001010101111011",
						 "000011001001011001101110",
						 "000011001001011101100001",
						 "000011001001100001010100",
						 "000011001001100101000111",
						 "000011001001101000111010",
						 "000011001001101100101101",
						 "000011001001110000100000",
						 "000011001001110100010011",
						 "000011001001111000000110",
						 "000011001001111011111001",
						 "000011001001111111101100",
						 "000011001010000011011111",
						 "000011001001001010100010",
						 "000011001001001110010100",
						 "000011001001010010000110",
						 "000011001001010101111000",
						 "000011001001011001101010",
						 "000011001001011101011100",
						 "000011001001100001001110",
						 "000011001001100101000000",
						 "000011001001101000110010",
						 "000011001001101100100100",
						 "000011001001110000010110",
						 "000011001001110100001000",
						 "000011001001110111111010",
						 "000011001001111011101100",
						 "000011001001111111011110",
						 "000011001010000011010000",
						 "000011001001001010100010",
						 "000011001001001110010100",
						 "000011001001010010000110",
						 "000011001001010101111000",
						 "000011001001011001101010",
						 "000011001001011101011100",
						 "000011001001100001001110",
						 "000011001001100101000000",
						 "000011001001101000110010",
						 "000011001001101100100100",
						 "000011001001110000010110",
						 "000011001001110100001000",
						 "000011001001110111111010",
						 "000011001001111011101100",
						 "000011001001111111011110",
						 "000011001010000011010000",
						 "000011001011101101100000",
						 "000011001011110001010010",
						 "000011001011110101000100",
						 "000011001011111000110110",
						 "000011001011111100101000",
						 "000011001100000000011010",
						 "000011001100000100001100",
						 "000011001100000111111110",
						 "000011001100001011110000",
						 "000011001100001111100010",
						 "000011001100010011010100",
						 "000011001100010111000110",
						 "000011001100011010111000",
						 "000011001100011110101010",
						 "000011001100100010011100",
						 "000011001100100110001110",
						 "000011001011101101100000",
						 "000011001011110001010010",
						 "000011001011110101000100",
						 "000011001011111000110110",
						 "000011001011111100101000",
						 "000011001100000000011010",
						 "000011001100000100001100",
						 "000011001100000111111110",
						 "000011001100001011110000",
						 "000011001100001111100010",
						 "000011001100010011010100",
						 "000011001100010111000110",
						 "000011001100011010111000",
						 "000011001100011110101010",
						 "000011001100100010011100",
						 "000011001100100110001110",
						 "000011001011101101100000",
						 "000011001011110001010010",
						 "000011001011110101000100",
						 "000011001011111000110110",
						 "000011001011111100101000",
						 "000011001100000000011010",
						 "000011001100000100001100",
						 "000011001100000111111110",
						 "000011001100001011110000",
						 "000011001100001111100010",
						 "000011001100010011010100",
						 "000011001100010111000110",
						 "000011001100011010111000",
						 "000011001100011110101010",
						 "000011001100100010011100",
						 "000011001100100110001110",
						 "000011001110010000011110",
						 "000011001110010100010000",
						 "000011001110011000000010",
						 "000011001110011011110100",
						 "000011001110011111100110",
						 "000011001110100011011000",
						 "000011001110100111001010",
						 "000011001110101010111100",
						 "000011001110101110101110",
						 "000011001110110010100000",
						 "000011001110110110010010",
						 "000011001110111010000100",
						 "000011001110111101110110",
						 "000011001111000001101000",
						 "000011001111000101011010",
						 "000011001111001001001100",
						 "000011001110010000011110",
						 "000011001110010100010000",
						 "000011001110011000000010",
						 "000011001110011011110100",
						 "000011001110011111100110",
						 "000011001110100011011000",
						 "000011001110100111001010",
						 "000011001110101010111100",
						 "000011001110101110101110",
						 "000011001110110010100000",
						 "000011001110110110010010",
						 "000011001110111010000100",
						 "000011001110111101110110",
						 "000011001111000001101000",
						 "000011001111000101011010",
						 "000011001111001001001100",
						 "000011001110010000011110",
						 "000011001110010100010000",
						 "000011001110011000000010",
						 "000011001110011011110100",
						 "000011001110011111100110",
						 "000011001110100011011000",
						 "000011001110100111001010",
						 "000011001110101010111100",
						 "000011001110101110101110",
						 "000011001110110010100000",
						 "000011001110110110010010",
						 "000011001110111010000100",
						 "000011001110111101110110",
						 "000011001111000001101000",
						 "000011001111000101011010",
						 "000011001111001001001100",
						 "000011010000110011011100",
						 "000011010000110111001101",
						 "000011010000111010111110",
						 "000011010000111110101111",
						 "000011010001000010100000",
						 "000011010001000110010001",
						 "000011010001001010000010",
						 "000011010001001101110011",
						 "000011010001010001100100",
						 "000011010001010101010101",
						 "000011010001011001000110",
						 "000011010001011100110111",
						 "000011010001100000101000",
						 "000011010001100100011001",
						 "000011010001101000001010",
						 "000011010001101011111011",
						 "000011010000110011011100",
						 "000011010000110111001101",
						 "000011010000111010111110",
						 "000011010000111110101111",
						 "000011010001000010100000",
						 "000011010001000110010001",
						 "000011010001001010000010",
						 "000011010001001101110011",
						 "000011010001010001100100",
						 "000011010001010101010101",
						 "000011010001011001000110",
						 "000011010001011100110111",
						 "000011010001100000101000",
						 "000011010001100100011001",
						 "000011010001101000001010",
						 "000011010001101011111011",
						 "000011010011010110011010",
						 "000011010011011010001011",
						 "000011010011011101111100",
						 "000011010011100001101101",
						 "000011010011100101011110",
						 "000011010011101001001111",
						 "000011010011101101000000",
						 "000011010011110000110001",
						 "000011010011110100100010",
						 "000011010011111000010011",
						 "000011010011111100000100",
						 "000011010011111111110101",
						 "000011010100000011100110",
						 "000011010100000111010111",
						 "000011010100001011001000",
						 "000011010100001110111001",
						 "000011010011010110011010",
						 "000011010011011010001011",
						 "000011010011011101111100",
						 "000011010011100001101101",
						 "000011010011100101011110",
						 "000011010011101001001111",
						 "000011010011101101000000",
						 "000011010011110000110001",
						 "000011010011110100100010",
						 "000011010011111000010011",
						 "000011010011111100000100",
						 "000011010011111111110101",
						 "000011010100000011100110",
						 "000011010100000111010111",
						 "000011010100001011001000",
						 "000011010100001110111001",
						 "000011010011010110011010",
						 "000011010011011010001011",
						 "000011010011011101111100",
						 "000011010011100001101101",
						 "000011010011100101011110",
						 "000011010011101001001111",
						 "000011010011101101000000",
						 "000011010011110000110001",
						 "000011010011110100100010",
						 "000011010011111000010011",
						 "000011010011111100000100",
						 "000011010011111111110101",
						 "000011010100000011100110",
						 "000011010100000111010111",
						 "000011010100001011001000",
						 "000011010100001110111001",
						 "000011010101111001011000",
						 "000011010101111101001001",
						 "000011010110000000111010",
						 "000011010110000100101011",
						 "000011010110001000011100",
						 "000011010110001100001101",
						 "000011010110001111111110",
						 "000011010110010011101111",
						 "000011010110010111100000",
						 "000011010110011011010001",
						 "000011010110011111000010",
						 "000011010110100010110011",
						 "000011010110100110100100",
						 "000011010110101010010101",
						 "000011010110101110000110",
						 "000011010110110001110111",
						 "000011010101111001011000",
						 "000011010101111101001001",
						 "000011010110000000111010",
						 "000011010110000100101011",
						 "000011010110001000011100",
						 "000011010110001100001101",
						 "000011010110001111111110",
						 "000011010110010011101111",
						 "000011010110010111100000",
						 "000011010110011011010001",
						 "000011010110011111000010",
						 "000011010110100010110011",
						 "000011010110100110100100",
						 "000011010110101010010101",
						 "000011010110101110000110",
						 "000011010110110001110111",
						 "000011010101111001011000",
						 "000011010101111101001001",
						 "000011010110000000111010",
						 "000011010110000100101011",
						 "000011010110001000011100",
						 "000011010110001100001101",
						 "000011010110001111111110",
						 "000011010110010011101111",
						 "000011010110010111100000",
						 "000011010110011011010001",
						 "000011010110011111000010",
						 "000011010110100010110011",
						 "000011010110100110100100",
						 "000011010110101010010101",
						 "000011010110101110000110",
						 "000011010110110001110111",
						 "000011011000011100010110",
						 "000011011000100000000110",
						 "000011011000100011110110",
						 "000011011000100111100110",
						 "000011011000101011010110",
						 "000011011000101111000110",
						 "000011011000110010110110",
						 "000011011000110110100110",
						 "000011011000111010010110",
						 "000011011000111110000110",
						 "000011011001000001110110",
						 "000011011001000101100110",
						 "000011011001001001010110",
						 "000011011001001101000110",
						 "000011011001010000110110",
						 "000011011001010100100110",
						 "000011011000011100010110",
						 "000011011000100000000110",
						 "000011011000100011110110",
						 "000011011000100111100110",
						 "000011011000101011010110",
						 "000011011000101111000110",
						 "000011011000110010110110",
						 "000011011000110110100110",
						 "000011011000111010010110",
						 "000011011000111110000110",
						 "000011011001000001110110",
						 "000011011001000101100110",
						 "000011011001001001010110",
						 "000011011001001101000110",
						 "000011011001010000110110",
						 "000011011001010100100110",
						 "000011011010111111010100",
						 "000011011011000011000100",
						 "000011011011000110110100",
						 "000011011011001010100100",
						 "000011011011001110010100",
						 "000011011011010010000100",
						 "000011011011010101110100",
						 "000011011011011001100100",
						 "000011011011011101010100",
						 "000011011011100001000100",
						 "000011011011100100110100",
						 "000011011011101000100100",
						 "000011011011101100010100",
						 "000011011011110000000100",
						 "000011011011110011110100",
						 "000011011011110111100100",
						 "000011011010111111010100",
						 "000011011011000011000100",
						 "000011011011000110110100",
						 "000011011011001010100100",
						 "000011011011001110010100",
						 "000011011011010010000100",
						 "000011011011010101110100",
						 "000011011011011001100100",
						 "000011011011011101010100",
						 "000011011011100001000100",
						 "000011011011100100110100",
						 "000011011011101000100100",
						 "000011011011101100010100",
						 "000011011011110000000100",
						 "000011011011110011110100",
						 "000011011011110111100100",
						 "000011011010111111010100",
						 "000011011011000011000100",
						 "000011011011000110110100",
						 "000011011011001010100100",
						 "000011011011001110010100",
						 "000011011011010010000100",
						 "000011011011010101110100",
						 "000011011011011001100100",
						 "000011011011011101010100",
						 "000011011011100001000100",
						 "000011011011100100110100",
						 "000011011011101000100100",
						 "000011011011101100010100",
						 "000011011011110000000100",
						 "000011011011110011110100",
						 "000011011011110111100100",
						 "000011011101100010010010",
						 "000011011101100110000010",
						 "000011011101101001110010",
						 "000011011101101101100010",
						 "000011011101110001010010",
						 "000011011101110101000010",
						 "000011011101111000110010",
						 "000011011101111100100010",
						 "000011011110000000010010",
						 "000011011110000100000010",
						 "000011011110000111110010",
						 "000011011110001011100010",
						 "000011011110001111010010",
						 "000011011110010011000010",
						 "000011011110010110110010",
						 "000011011110011010100010",
						 "000011011101100010010010",
						 "000011011101100110000010",
						 "000011011101101001110010",
						 "000011011101101101100010",
						 "000011011101110001010010",
						 "000011011101110101000010",
						 "000011011101111000110010",
						 "000011011101111100100010",
						 "000011011110000000010010",
						 "000011011110000100000010",
						 "000011011110000111110010",
						 "000011011110001011100010",
						 "000011011110001111010010",
						 "000011011110010011000010",
						 "000011011110010110110010",
						 "000011011110011010100010",
						 "000011011101100010010010",
						 "000011011101100110000001",
						 "000011011101101001110000",
						 "000011011101101101011111",
						 "000011011101110001001110",
						 "000011011101110100111101",
						 "000011011101111000101100",
						 "000011011101111100011011",
						 "000011011110000000001010",
						 "000011011110000011111001",
						 "000011011110000111101000",
						 "000011011110001011010111",
						 "000011011110001111000110",
						 "000011011110010010110101",
						 "000011011110010110100100",
						 "000011011110011010010011",
						 "000011100000000101010000",
						 "000011100000001000111111",
						 "000011100000001100101110",
						 "000011100000010000011101",
						 "000011100000010100001100",
						 "000011100000010111111011",
						 "000011100000011011101010",
						 "000011100000011111011001",
						 "000011100000100011001000",
						 "000011100000100110110111",
						 "000011100000101010100110",
						 "000011100000101110010101",
						 "000011100000110010000100",
						 "000011100000110101110011",
						 "000011100000111001100010",
						 "000011100000111101010001",
						 "000011100000000101010000",
						 "000011100000001000111111",
						 "000011100000001100101110",
						 "000011100000010000011101",
						 "000011100000010100001100",
						 "000011100000010111111011",
						 "000011100000011011101010",
						 "000011100000011111011001",
						 "000011100000100011001000",
						 "000011100000100110110111",
						 "000011100000101010100110",
						 "000011100000101110010101",
						 "000011100000110010000100",
						 "000011100000110101110011",
						 "000011100000111001100010",
						 "000011100000111101010001",
						 "000011100000000101010000",
						 "000011100000001000111111",
						 "000011100000001100101110",
						 "000011100000010000011101",
						 "000011100000010100001100",
						 "000011100000010111111011",
						 "000011100000011011101010",
						 "000011100000011111011001",
						 "000011100000100011001000",
						 "000011100000100110110111",
						 "000011100000101010100110",
						 "000011100000101110010101",
						 "000011100000110010000100",
						 "000011100000110101110011",
						 "000011100000111001100010",
						 "000011100000111101010001",
						 "000011100010101000001110",
						 "000011100010101011111101",
						 "000011100010101111101100",
						 "000011100010110011011011",
						 "000011100010110111001010",
						 "000011100010111010111001",
						 "000011100010111110101000",
						 "000011100011000010010111",
						 "000011100011000110000110",
						 "000011100011001001110101",
						 "000011100011001101100100",
						 "000011100011010001010011",
						 "000011100011010101000010",
						 "000011100011011000110001",
						 "000011100011011100100000",
						 "000011100011100000001111",
						 "000011100010101000001110",
						 "000011100010101011111101",
						 "000011100010101111101100",
						 "000011100010110011011011",
						 "000011100010110111001010",
						 "000011100010111010111001",
						 "000011100010111110101000",
						 "000011100011000010010111",
						 "000011100011000110000110",
						 "000011100011001001110101",
						 "000011100011001101100100",
						 "000011100011010001010011",
						 "000011100011010101000010",
						 "000011100011011000110001",
						 "000011100011011100100000",
						 "000011100011100000001111",
						 "000011100101001011001100",
						 "000011100101001110111011",
						 "000011100101010010101010",
						 "000011100101010110011001",
						 "000011100101011010001000",
						 "000011100101011101110111",
						 "000011100101100001100110",
						 "000011100101100101010101",
						 "000011100101101001000100",
						 "000011100101101100110011",
						 "000011100101110000100010",
						 "000011100101110100010001",
						 "000011100101111000000000",
						 "000011100101111011101111",
						 "000011100101111111011110",
						 "000011100110000011001101",
						 "000011100101001011001100",
						 "000011100101001110111011",
						 "000011100101010010101010",
						 "000011100101010110011001",
						 "000011100101011010001000",
						 "000011100101011101110111",
						 "000011100101100001100110",
						 "000011100101100101010101",
						 "000011100101101001000100",
						 "000011100101101100110011",
						 "000011100101110000100010",
						 "000011100101110100010001",
						 "000011100101111000000000",
						 "000011100101111011101111",
						 "000011100101111111011110",
						 "000011100110000011001101",
						 "000011100101001011001100",
						 "000011100101001110111010",
						 "000011100101010010101000",
						 "000011100101010110010110",
						 "000011100101011010000100",
						 "000011100101011101110010",
						 "000011100101100001100000",
						 "000011100101100101001110",
						 "000011100101101000111100",
						 "000011100101101100101010",
						 "000011100101110000011000",
						 "000011100101110100000110",
						 "000011100101110111110100",
						 "000011100101111011100010",
						 "000011100101111111010000",
						 "000011100110000010111110",
						 "000011100111101110001010",
						 "000011100111110001111000",
						 "000011100111110101100110",
						 "000011100111111001010100",
						 "000011100111111101000010",
						 "000011101000000000110000",
						 "000011101000000100011110",
						 "000011101000001000001100",
						 "000011101000001011111010",
						 "000011101000001111101000",
						 "000011101000010011010110",
						 "000011101000010111000100",
						 "000011101000011010110010",
						 "000011101000011110100000",
						 "000011101000100010001110",
						 "000011101000100101111100",
						 "000011100111101110001010",
						 "000011100111110001111000",
						 "000011100111110101100110",
						 "000011100111111001010100",
						 "000011100111111101000010",
						 "000011101000000000110000",
						 "000011101000000100011110",
						 "000011101000001000001100",
						 "000011101000001011111010",
						 "000011101000001111101000",
						 "000011101000010011010110",
						 "000011101000010111000100",
						 "000011101000011010110010",
						 "000011101000011110100000",
						 "000011101000100010001110",
						 "000011101000100101111100",
						 "000011100111101110001010",
						 "000011100111110001111000",
						 "000011100111110101100110",
						 "000011100111111001010100",
						 "000011100111111101000010",
						 "000011101000000000110000",
						 "000011101000000100011110",
						 "000011101000001000001100",
						 "000011101000001011111010",
						 "000011101000001111101000",
						 "000011101000010011010110",
						 "000011101000010111000100",
						 "000011101000011010110010",
						 "000011101000011110100000",
						 "000011101000100010001110",
						 "000011101000100101111100",
						 "000011101010010001001000",
						 "000011101010010100110110",
						 "000011101010011000100100",
						 "000011101010011100010010",
						 "000011101010100000000000",
						 "000011101010100011101110",
						 "000011101010100111011100",
						 "000011101010101011001010",
						 "000011101010101110111000",
						 "000011101010110010100110",
						 "000011101010110110010100",
						 "000011101010111010000010",
						 "000011101010111101110000",
						 "000011101011000001011110",
						 "000011101011000101001100",
						 "000011101011001000111010",
						 "000011101010010001001000",
						 "000011101010010100110110",
						 "000011101010011000100100",
						 "000011101010011100010010",
						 "000011101010100000000000",
						 "000011101010100011101110",
						 "000011101010100111011100",
						 "000011101010101011001010",
						 "000011101010101110111000",
						 "000011101010110010100110",
						 "000011101010110110010100",
						 "000011101010111010000010",
						 "000011101010111101110000",
						 "000011101011000001011110",
						 "000011101011000101001100",
						 "000011101011001000111010",
						 "000011101100110100000110",
						 "000011101100110111110100",
						 "000011101100111011100010",
						 "000011101100111111010000",
						 "000011101101000010111110",
						 "000011101101000110101100",
						 "000011101101001010011010",
						 "000011101101001110001000",
						 "000011101101010001110110",
						 "000011101101010101100100",
						 "000011101101011001010010",
						 "000011101101011101000000",
						 "000011101101100000101110",
						 "000011101101100100011100",
						 "000011101101101000001010",
						 "000011101101101011111000",
						 "000011101100110100000110",
						 "000011101100110111110011",
						 "000011101100111011100000",
						 "000011101100111111001101",
						 "000011101101000010111010",
						 "000011101101000110100111",
						 "000011101101001010010100",
						 "000011101101001110000001",
						 "000011101101010001101110",
						 "000011101101010101011011",
						 "000011101101011001001000",
						 "000011101101011100110101",
						 "000011101101100000100010",
						 "000011101101100100001111",
						 "000011101101100111111100",
						 "000011101101101011101001",
						 "000011101100110100000110",
						 "000011101100110111110011",
						 "000011101100111011100000",
						 "000011101100111111001101",
						 "000011101101000010111010",
						 "000011101101000110100111",
						 "000011101101001010010100",
						 "000011101101001110000001",
						 "000011101101010001101110",
						 "000011101101010101011011",
						 "000011101101011001001000",
						 "000011101101011100110101",
						 "000011101101100000100010",
						 "000011101101100100001111",
						 "000011101101100111111100",
						 "000011101101101011101001",
						 "000011101111010111000100",
						 "000011101111011010110001",
						 "000011101111011110011110",
						 "000011101111100010001011",
						 "000011101111100101111000",
						 "000011101111101001100101",
						 "000011101111101101010010",
						 "000011101111110000111111",
						 "000011101111110100101100",
						 "000011101111111000011001",
						 "000011101111111100000110",
						 "000011101111111111110011",
						 "000011110000000011100000",
						 "000011110000000111001101",
						 "000011110000001010111010",
						 "000011110000001110100111",
						 "000011101111010111000100",
						 "000011101111011010110001",
						 "000011101111011110011110",
						 "000011101111100010001011",
						 "000011101111100101111000",
						 "000011101111101001100101",
						 "000011101111101101010010",
						 "000011101111110000111111",
						 "000011101111110100101100",
						 "000011101111111000011001",
						 "000011101111111100000110",
						 "000011101111111111110011",
						 "000011110000000011100000",
						 "000011110000000111001101",
						 "000011110000001010111010",
						 "000011110000001110100111",
						 "000011101111010111000100",
						 "000011101111011010110001",
						 "000011101111011110011110",
						 "000011101111100010001011",
						 "000011101111100101111000",
						 "000011101111101001100101",
						 "000011101111101101010010",
						 "000011101111110000111111",
						 "000011101111110100101100",
						 "000011101111111000011001",
						 "000011101111111100000110",
						 "000011101111111111110011",
						 "000011110000000011100000",
						 "000011110000000111001101",
						 "000011110000001010111010",
						 "000011110000001110100111",
						 "000011110001111010000010",
						 "000011110001111101101111",
						 "000011110010000001011100",
						 "000011110010000101001001",
						 "000011110010001000110110",
						 "000011110010001100100011",
						 "000011110010010000010000",
						 "000011110010010011111101",
						 "000011110010010111101010",
						 "000011110010011011010111",
						 "000011110010011111000100",
						 "000011110010100010110001",
						 "000011110010100110011110",
						 "000011110010101010001011",
						 "000011110010101101111000",
						 "000011110010110001100101",
						 "000011110001111010000010",
						 "000011110001111101101111",
						 "000011110010000001011100",
						 "000011110010000101001001",
						 "000011110010001000110110",
						 "000011110010001100100011",
						 "000011110010010000010000",
						 "000011110010010011111101",
						 "000011110010010111101010",
						 "000011110010011011010111",
						 "000011110010011111000100",
						 "000011110010100010110001",
						 "000011110010100110011110",
						 "000011110010101010001011",
						 "000011110010101101111000",
						 "000011110010110001100101",
						 "000011110001111010000010",
						 "000011110001111101101110",
						 "000011110010000001011010",
						 "000011110010000101000110",
						 "000011110010001000110010",
						 "000011110010001100011110",
						 "000011110010010000001010",
						 "000011110010010011110110",
						 "000011110010010111100010",
						 "000011110010011011001110",
						 "000011110010011110111010",
						 "000011110010100010100110",
						 "000011110010100110010010",
						 "000011110010101001111110",
						 "000011110010101101101010",
						 "000011110010110001010110",
						 "000011110100011101000000",
						 "000011110100100000101100",
						 "000011110100100100011000",
						 "000011110100101000000100",
						 "000011110100101011110000",
						 "000011110100101111011100",
						 "000011110100110011001000",
						 "000011110100110110110100",
						 "000011110100111010100000",
						 "000011110100111110001100",
						 "000011110101000001111000",
						 "000011110101000101100100",
						 "000011110101001001010000",
						 "000011110101001100111100",
						 "000011110101010000101000",
						 "000011110101010100010100",
						 "000011110100011101000000",
						 "000011110100100000101100",
						 "000011110100100100011000",
						 "000011110100101000000100",
						 "000011110100101011110000",
						 "000011110100101111011100",
						 "000011110100110011001000",
						 "000011110100110110110100",
						 "000011110100111010100000",
						 "000011110100111110001100",
						 "000011110101000001111000",
						 "000011110101000101100100",
						 "000011110101001001010000",
						 "000011110101001100111100",
						 "000011110101010000101000",
						 "000011110101010100010100",
						 "000011110110111111111110",
						 "000011110111000011101010",
						 "000011110111000111010110",
						 "000011110111001011000010",
						 "000011110111001110101110",
						 "000011110111010010011010",
						 "000011110111010110000110",
						 "000011110111011001110010",
						 "000011110111011101011110",
						 "000011110111100001001010",
						 "000011110111100100110110",
						 "000011110111101000100010",
						 "000011110111101100001110",
						 "000011110111101111111010",
						 "000011110111110011100110",
						 "000011110111110111010010",
						 "000011110110111111111110",
						 "000011110111000011101010",
						 "000011110111000111010110",
						 "000011110111001011000010",
						 "000011110111001110101110",
						 "000011110111010010011010",
						 "000011110111010110000110",
						 "000011110111011001110010",
						 "000011110111011101011110",
						 "000011110111100001001010",
						 "000011110111100100110110",
						 "000011110111101000100010",
						 "000011110111101100001110",
						 "000011110111101111111010",
						 "000011110111110011100110",
						 "000011110111110111010010",
						 "000011110110111111111110",
						 "000011110111000011101010",
						 "000011110111000111010110",
						 "000011110111001011000010",
						 "000011110111001110101110",
						 "000011110111010010011010",
						 "000011110111010110000110",
						 "000011110111011001110010",
						 "000011110111011101011110",
						 "000011110111100001001010",
						 "000011110111100100110110",
						 "000011110111101000100010",
						 "000011110111101100001110",
						 "000011110111101111111010",
						 "000011110111110011100110",
						 "000011110111110111010010",
						 "000011111001100010111100",
						 "000011111001100110101000",
						 "000011111001101010010100",
						 "000011111001101110000000",
						 "000011111001110001101100",
						 "000011111001110101011000",
						 "000011111001111001000100",
						 "000011111001111100110000",
						 "000011111010000000011100",
						 "000011111010000100001000",
						 "000011111010000111110100",
						 "000011111010001011100000",
						 "000011111010001111001100",
						 "000011111010010010111000",
						 "000011111010010110100100",
						 "000011111010011010010000",
						 "000011111001100010111100",
						 "000011111001100110100111",
						 "000011111001101010010010",
						 "000011111001101101111101",
						 "000011111001110001101000",
						 "000011111001110101010011",
						 "000011111001111000111110",
						 "000011111001111100101001",
						 "000011111010000000010100",
						 "000011111010000011111111",
						 "000011111010000111101010",
						 "000011111010001011010101",
						 "000011111010001111000000",
						 "000011111010010010101011",
						 "000011111010010110010110",
						 "000011111010011010000001",
						 "000011111001100010111100",
						 "000011111001100110100111",
						 "000011111001101010010010",
						 "000011111001101101111101",
						 "000011111001110001101000",
						 "000011111001110101010011",
						 "000011111001111000111110",
						 "000011111001111100101001",
						 "000011111010000000010100",
						 "000011111010000011111111",
						 "000011111010000111101010",
						 "000011111010001011010101",
						 "000011111010001111000000",
						 "000011111010010010101011",
						 "000011111010010110010110",
						 "000011111010011010000001",
						 "000011111100000101111010",
						 "000011111100001001100101",
						 "000011111100001101010000",
						 "000011111100010000111011",
						 "000011111100010100100110",
						 "000011111100011000010001",
						 "000011111100011011111100",
						 "000011111100011111100111",
						 "000011111100100011010010",
						 "000011111100100110111101",
						 "000011111100101010101000",
						 "000011111100101110010011",
						 "000011111100110001111110",
						 "000011111100110101101001",
						 "000011111100111001010100",
						 "000011111100111100111111",
						 "000011111100000101111010",
						 "000011111100001001100101",
						 "000011111100001101010000",
						 "000011111100010000111011",
						 "000011111100010100100110",
						 "000011111100011000010001",
						 "000011111100011011111100",
						 "000011111100011111100111",
						 "000011111100100011010010",
						 "000011111100100110111101",
						 "000011111100101010101000",
						 "000011111100101110010011",
						 "000011111100110001111110",
						 "000011111100110101101001",
						 "000011111100111001010100",
						 "000011111100111100111111",
						 "000011111100000101111010",
						 "000011111100001001100101",
						 "000011111100001101010000",
						 "000011111100010000111011",
						 "000011111100010100100110",
						 "000011111100011000010001",
						 "000011111100011011111100",
						 "000011111100011111100111",
						 "000011111100100011010010",
						 "000011111100100110111101",
						 "000011111100101010101000",
						 "000011111100101110010011",
						 "000011111100110001111110",
						 "000011111100110101101001",
						 "000011111100111001010100",
						 "000011111100111100111111",
						 "000011111110101000111000",
						 "000011111110101100100011",
						 "000011111110110000001110",
						 "000011111110110011111001",
						 "000011111110110111100100",
						 "000011111110111011001111",
						 "000011111110111110111010",
						 "000011111111000010100101",
						 "000011111111000110010000",
						 "000011111111001001111011",
						 "000011111111001101100110",
						 "000011111111010001010001",
						 "000011111111010100111100",
						 "000011111111011000100111",
						 "000011111111011100010010",
						 "000011111111011111111101",
						 "000011111110101000111000",
						 "000011111110101100100010",
						 "000011111110110000001100",
						 "000011111110110011110110",
						 "000011111110110111100000",
						 "000011111110111011001010",
						 "000011111110111110110100",
						 "000011111111000010011110",
						 "000011111111000110001000",
						 "000011111111001001110010",
						 "000011111111001101011100",
						 "000011111111010001000110",
						 "000011111111010100110000",
						 "000011111111011000011010",
						 "000011111111011100000100",
						 "000011111111011111101110",
						 "000011111110101000111000",
						 "000011111110101100100010",
						 "000011111110110000001100",
						 "000011111110110011110110",
						 "000011111110110111100000",
						 "000011111110111011001010",
						 "000011111110111110110100",
						 "000011111111000010011110",
						 "000011111111000110001000",
						 "000011111111001001110010",
						 "000011111111001101011100",
						 "000011111111010001000110",
						 "000011111111010100110000",
						 "000011111111011000011010",
						 "000011111111011100000100",
						 "000011111111011111101110",
						 "000100000001001011110110",
						 "000100000001001111100000",
						 "000100000001010011001010",
						 "000100000001010110110100",
						 "000100000001011010011110",
						 "000100000001011110001000",
						 "000100000001100001110010",
						 "000100000001100101011100",
						 "000100000001101001000110",
						 "000100000001101100110000",
						 "000100000001110000011010",
						 "000100000001110100000100",
						 "000100000001110111101110",
						 "000100000001111011011000",
						 "000100000001111111000010",
						 "000100000010000010101100",
						 "000100000001001011110110",
						 "000100000001001111100000",
						 "000100000001010011001010",
						 "000100000001010110110100",
						 "000100000001011010011110",
						 "000100000001011110001000",
						 "000100000001100001110010",
						 "000100000001100101011100",
						 "000100000001101001000110",
						 "000100000001101100110000",
						 "000100000001110000011010",
						 "000100000001110100000100",
						 "000100000001110111101110",
						 "000100000001111011011000",
						 "000100000001111111000010",
						 "000100000010000010101100",
						 "000100000011101110110100",
						 "000100000011110010011110",
						 "000100000011110110001000",
						 "000100000011111001110010",
						 "000100000011111101011100",
						 "000100000100000001000110",
						 "000100000100000100110000",
						 "000100000100001000011010",
						 "000100000100001100000100",
						 "000100000100001111101110",
						 "000100000100010011011000",
						 "000100000100010111000010",
						 "000100000100011010101100",
						 "000100000100011110010110",
						 "000100000100100010000000",
						 "000100000100100101101010",
						 "000100000011101110110100",
						 "000100000011110010011110",
						 "000100000011110110001000",
						 "000100000011111001110010",
						 "000100000011111101011100",
						 "000100000100000001000110",
						 "000100000100000100110000",
						 "000100000100001000011010",
						 "000100000100001100000100",
						 "000100000100001111101110",
						 "000100000100010011011000",
						 "000100000100010111000010",
						 "000100000100011010101100",
						 "000100000100011110010110",
						 "000100000100100010000000",
						 "000100000100100101101010",
						 "000100000011101110110100",
						 "000100000011110010011110",
						 "000100000011110110001000",
						 "000100000011111001110010",
						 "000100000011111101011100",
						 "000100000100000001000110",
						 "000100000100000100110000",
						 "000100000100001000011010",
						 "000100000100001100000100",
						 "000100000100001111101110",
						 "000100000100010011011000",
						 "000100000100010111000010",
						 "000100000100011010101100",
						 "000100000100011110010110",
						 "000100000100100010000000",
						 "000100000100100101101010",
						 "000100000110010001110010",
						 "000100000110010101011011",
						 "000100000110011001000100",
						 "000100000110011100101101",
						 "000100000110100000010110",
						 "000100000110100011111111",
						 "000100000110100111101000",
						 "000100000110101011010001",
						 "000100000110101110111010",
						 "000100000110110010100011",
						 "000100000110110110001100",
						 "000100000110111001110101",
						 "000100000110111101011110",
						 "000100000111000001000111",
						 "000100000111000100110000",
						 "000100000111001000011001",
						 "000100000110010001110010",
						 "000100000110010101011011",
						 "000100000110011001000100",
						 "000100000110011100101101",
						 "000100000110100000010110",
						 "000100000110100011111111",
						 "000100000110100111101000",
						 "000100000110101011010001",
						 "000100000110101110111010",
						 "000100000110110010100011",
						 "000100000110110110001100",
						 "000100000110111001110101",
						 "000100000110111101011110",
						 "000100000111000001000111",
						 "000100000111000100110000",
						 "000100000111001000011001",
						 "000100000110010001110010",
						 "000100000110010101011011",
						 "000100000110011001000100",
						 "000100000110011100101101",
						 "000100000110100000010110",
						 "000100000110100011111111",
						 "000100000110100111101000",
						 "000100000110101011010001",
						 "000100000110101110111010",
						 "000100000110110010100011",
						 "000100000110110110001100",
						 "000100000110111001110101",
						 "000100000110111101011110",
						 "000100000111000001000111",
						 "000100000111000100110000",
						 "000100000111001000011001",
						 "000100001000110100110000",
						 "000100001000111000011001",
						 "000100001000111100000010",
						 "000100001000111111101011",
						 "000100001001000011010100",
						 "000100001001000110111101",
						 "000100001001001010100110",
						 "000100001001001110001111",
						 "000100001001010001111000",
						 "000100001001010101100001",
						 "000100001001011001001010",
						 "000100001001011100110011",
						 "000100001001100000011100",
						 "000100001001100100000101",
						 "000100001001100111101110",
						 "000100001001101011010111",
						 "000100001000110100110000",
						 "000100001000111000011001",
						 "000100001000111100000010",
						 "000100001000111111101011",
						 "000100001001000011010100",
						 "000100001001000110111101",
						 "000100001001001010100110",
						 "000100001001001110001111",
						 "000100001001010001111000",
						 "000100001001010101100001",
						 "000100001001011001001010",
						 "000100001001011100110011",
						 "000100001001100000011100",
						 "000100001001100100000101",
						 "000100001001100111101110",
						 "000100001001101011010111",
						 "000100001000110100110000",
						 "000100001000111000011001",
						 "000100001000111100000010",
						 "000100001000111111101011",
						 "000100001001000011010100",
						 "000100001001000110111101",
						 "000100001001001010100110",
						 "000100001001001110001111",
						 "000100001001010001111000",
						 "000100001001010101100001",
						 "000100001001011001001010",
						 "000100001001011100110011",
						 "000100001001100000011100",
						 "000100001001100100000101",
						 "000100001001100111101110",
						 "000100001001101011010111",
						 "000100001011010111101110",
						 "000100001011011011010110",
						 "000100001011011110111110",
						 "000100001011100010100110",
						 "000100001011100110001110",
						 "000100001011101001110110",
						 "000100001011101101011110",
						 "000100001011110001000110",
						 "000100001011110100101110",
						 "000100001011111000010110",
						 "000100001011111011111110",
						 "000100001011111111100110",
						 "000100001100000011001110",
						 "000100001100000110110110",
						 "000100001100001010011110",
						 "000100001100001110000110",
						 "000100001011010111101110",
						 "000100001011011011010110",
						 "000100001011011110111110",
						 "000100001011100010100110",
						 "000100001011100110001110",
						 "000100001011101001110110",
						 "000100001011101101011110",
						 "000100001011110001000110",
						 "000100001011110100101110",
						 "000100001011111000010110",
						 "000100001011111011111110",
						 "000100001011111111100110",
						 "000100001100000011001110",
						 "000100001100000110110110",
						 "000100001100001010011110",
						 "000100001100001110000110",
						 "000100001011010111101110",
						 "000100001011011011010110",
						 "000100001011011110111110",
						 "000100001011100010100110",
						 "000100001011100110001110",
						 "000100001011101001110110",
						 "000100001011101101011110",
						 "000100001011110001000110",
						 "000100001011110100101110",
						 "000100001011111000010110",
						 "000100001011111011111110",
						 "000100001011111111100110",
						 "000100001100000011001110",
						 "000100001100000110110110",
						 "000100001100001010011110",
						 "000100001100001110000110",
						 "000100001101111010101100",
						 "000100001101111110010100",
						 "000100001110000001111100",
						 "000100001110000101100100",
						 "000100001110001001001100",
						 "000100001110001100110100",
						 "000100001110010000011100",
						 "000100001110010100000100",
						 "000100001110010111101100",
						 "000100001110011011010100",
						 "000100001110011110111100",
						 "000100001110100010100100",
						 "000100001110100110001100",
						 "000100001110101001110100",
						 "000100001110101101011100",
						 "000100001110110001000100",
						 "000100001101111010101100",
						 "000100001101111110010100",
						 "000100001110000001111100",
						 "000100001110000101100100",
						 "000100001110001001001100",
						 "000100001110001100110100",
						 "000100001110010000011100",
						 "000100001110010100000100",
						 "000100001110010111101100",
						 "000100001110011011010100",
						 "000100001110011110111100",
						 "000100001110100010100100",
						 "000100001110100110001100",
						 "000100001110101001110100",
						 "000100001110101101011100",
						 "000100001110110001000100",
						 "000100010000011101101010",
						 "000100010000100001010010",
						 "000100010000100100111010",
						 "000100010000101000100010",
						 "000100010000101100001010",
						 "000100010000101111110010",
						 "000100010000110011011010",
						 "000100010000110111000010",
						 "000100010000111010101010",
						 "000100010000111110010010",
						 "000100010001000001111010",
						 "000100010001000101100010",
						 "000100010001001001001010",
						 "000100010001001100110010",
						 "000100010001010000011010",
						 "000100010001010100000010",
						 "000100010000011101101010",
						 "000100010000100001010001",
						 "000100010000100100111000",
						 "000100010000101000011111",
						 "000100010000101100000110",
						 "000100010000101111101101",
						 "000100010000110011010100",
						 "000100010000110110111011",
						 "000100010000111010100010",
						 "000100010000111110001001",
						 "000100010001000001110000",
						 "000100010001000101010111",
						 "000100010001001000111110",
						 "000100010001001100100101",
						 "000100010001010000001100",
						 "000100010001010011110011",
						 "000100010000011101101010",
						 "000100010000100001010001",
						 "000100010000100100111000",
						 "000100010000101000011111",
						 "000100010000101100000110",
						 "000100010000101111101101",
						 "000100010000110011010100",
						 "000100010000110110111011",
						 "000100010000111010100010",
						 "000100010000111110001001",
						 "000100010001000001110000",
						 "000100010001000101010111",
						 "000100010001001000111110",
						 "000100010001001100100101",
						 "000100010001010000001100",
						 "000100010001010011110011",
						 "000100010011000000101000",
						 "000100010011000100001111",
						 "000100010011000111110110",
						 "000100010011001011011101",
						 "000100010011001111000100",
						 "000100010011010010101011",
						 "000100010011010110010010",
						 "000100010011011001111001",
						 "000100010011011101100000",
						 "000100010011100001000111",
						 "000100010011100100101110",
						 "000100010011101000010101",
						 "000100010011101011111100",
						 "000100010011101111100011",
						 "000100010011110011001010",
						 "000100010011110110110001",
						 "000100010011000000101000",
						 "000100010011000100001111",
						 "000100010011000111110110",
						 "000100010011001011011101",
						 "000100010011001111000100",
						 "000100010011010010101011",
						 "000100010011010110010010",
						 "000100010011011001111001",
						 "000100010011011101100000",
						 "000100010011100001000111",
						 "000100010011100100101110",
						 "000100010011101000010101",
						 "000100010011101011111100",
						 "000100010011101111100011",
						 "000100010011110011001010",
						 "000100010011110110110001",
						 "000100010011000000101000",
						 "000100010011000100001111",
						 "000100010011000111110110",
						 "000100010011001011011101",
						 "000100010011001111000100",
						 "000100010011010010101011",
						 "000100010011010110010010",
						 "000100010011011001111001",
						 "000100010011011101100000",
						 "000100010011100001000111",
						 "000100010011100100101110",
						 "000100010011101000010101",
						 "000100010011101011111100",
						 "000100010011101111100011",
						 "000100010011110011001010",
						 "000100010011110110110001",
						 "000100010101100011100110",
						 "000100010101100111001101",
						 "000100010101101010110100",
						 "000100010101101110011011",
						 "000100010101110010000010",
						 "000100010101110101101001",
						 "000100010101111001010000",
						 "000100010101111100110111",
						 "000100010110000000011110",
						 "000100010110000100000101",
						 "000100010110000111101100",
						 "000100010110001011010011",
						 "000100010110001110111010",
						 "000100010110010010100001",
						 "000100010110010110001000",
						 "000100010110011001101111",
						 "000100010101100011100110",
						 "000100010101100111001100",
						 "000100010101101010110010",
						 "000100010101101110011000",
						 "000100010101110001111110",
						 "000100010101110101100100",
						 "000100010101111001001010",
						 "000100010101111100110000",
						 "000100010110000000010110",
						 "000100010110000011111100",
						 "000100010110000111100010",
						 "000100010110001011001000",
						 "000100010110001110101110",
						 "000100010110010010010100",
						 "000100010110010101111010",
						 "000100010110011001100000",
						 "000100010101100011100110",
						 "000100010101100111001100",
						 "000100010101101010110010",
						 "000100010101101110011000",
						 "000100010101110001111110",
						 "000100010101110101100100",
						 "000100010101111001001010",
						 "000100010101111100110000",
						 "000100010110000000010110",
						 "000100010110000011111100",
						 "000100010110000111100010",
						 "000100010110001011001000",
						 "000100010110001110101110",
						 "000100010110010010010100",
						 "000100010110010101111010",
						 "000100010110011001100000",
						 "000100011000000110100100",
						 "000100011000001010001010",
						 "000100011000001101110000",
						 "000100011000010001010110",
						 "000100011000010100111100",
						 "000100011000011000100010",
						 "000100011000011100001000",
						 "000100011000011111101110",
						 "000100011000100011010100",
						 "000100011000100110111010",
						 "000100011000101010100000",
						 "000100011000101110000110",
						 "000100011000110001101100",
						 "000100011000110101010010",
						 "000100011000111000111000",
						 "000100011000111100011110",
						 "000100011000000110100100",
						 "000100011000001010001010",
						 "000100011000001101110000",
						 "000100011000010001010110",
						 "000100011000010100111100",
						 "000100011000011000100010",
						 "000100011000011100001000",
						 "000100011000011111101110",
						 "000100011000100011010100",
						 "000100011000100110111010",
						 "000100011000101010100000",
						 "000100011000101110000110",
						 "000100011000110001101100",
						 "000100011000110101010010",
						 "000100011000111000111000",
						 "000100011000111100011110",
						 "000100011000000110100100",
						 "000100011000001010001010",
						 "000100011000001101110000",
						 "000100011000010001010110",
						 "000100011000010100111100",
						 "000100011000011000100010",
						 "000100011000011100001000",
						 "000100011000011111101110",
						 "000100011000100011010100",
						 "000100011000100110111010",
						 "000100011000101010100000",
						 "000100011000101110000110",
						 "000100011000110001101100",
						 "000100011000110101010010",
						 "000100011000111000111000",
						 "000100011000111100011110",
						 "000100011010101001100010",
						 "000100011010101101001000",
						 "000100011010110000101110",
						 "000100011010110100010100",
						 "000100011010110111111010",
						 "000100011010111011100000",
						 "000100011010111111000110",
						 "000100011011000010101100",
						 "000100011011000110010010",
						 "000100011011001001111000",
						 "000100011011001101011110",
						 "000100011011010001000100",
						 "000100011011010100101010",
						 "000100011011011000010000",
						 "000100011011011011110110",
						 "000100011011011111011100",
						 "000100011010101001100010",
						 "000100011010101101000111",
						 "000100011010110000101100",
						 "000100011010110100010001",
						 "000100011010110111110110",
						 "000100011010111011011011",
						 "000100011010111111000000",
						 "000100011011000010100101",
						 "000100011011000110001010",
						 "000100011011001001101111",
						 "000100011011001101010100",
						 "000100011011010000111001",
						 "000100011011010100011110",
						 "000100011011011000000011",
						 "000100011011011011101000",
						 "000100011011011111001101",
						 "000100011010101001100010",
						 "000100011010101101000111",
						 "000100011010110000101100",
						 "000100011010110100010001",
						 "000100011010110111110110",
						 "000100011010111011011011",
						 "000100011010111111000000",
						 "000100011011000010100101",
						 "000100011011000110001010",
						 "000100011011001001101111",
						 "000100011011001101010100",
						 "000100011011010000111001",
						 "000100011011010100011110",
						 "000100011011011000000011",
						 "000100011011011011101000",
						 "000100011011011111001101",
						 "000100011101001100100000",
						 "000100011101010000000101",
						 "000100011101010011101010",
						 "000100011101010111001111",
						 "000100011101011010110100",
						 "000100011101011110011001",
						 "000100011101100001111110",
						 "000100011101100101100011",
						 "000100011101101001001000",
						 "000100011101101100101101",
						 "000100011101110000010010",
						 "000100011101110011110111",
						 "000100011101110111011100",
						 "000100011101111011000001",
						 "000100011101111110100110",
						 "000100011110000010001011",
						 "000100011101001100100000",
						 "000100011101010000000101",
						 "000100011101010011101010",
						 "000100011101010111001111",
						 "000100011101011010110100",
						 "000100011101011110011001",
						 "000100011101100001111110",
						 "000100011101100101100011",
						 "000100011101101001001000",
						 "000100011101101100101101",
						 "000100011101110000010010",
						 "000100011101110011110111",
						 "000100011101110111011100",
						 "000100011101111011000001",
						 "000100011101111110100110",
						 "000100011110000010001011",
						 "000100011111101111011110",
						 "000100011111110011000011",
						 "000100011111110110101000",
						 "000100011111111010001101",
						 "000100011111111101110010",
						 "000100100000000001010111",
						 "000100100000000100111100",
						 "000100100000001000100001",
						 "000100100000001100000110",
						 "000100100000001111101011",
						 "000100100000010011010000",
						 "000100100000010110110101",
						 "000100100000011010011010",
						 "000100100000011101111111",
						 "000100100000100001100100",
						 "000100100000100101001001",
						 "000100011111101111011110",
						 "000100011111110011000011",
						 "000100011111110110101000",
						 "000100011111111010001101",
						 "000100011111111101110010",
						 "000100100000000001010111",
						 "000100100000000100111100",
						 "000100100000001000100001",
						 "000100100000001100000110",
						 "000100100000001111101011",
						 "000100100000010011010000",
						 "000100100000010110110101",
						 "000100100000011010011010",
						 "000100100000011101111111",
						 "000100100000100001100100",
						 "000100100000100101001001",
						 "000100011111101111011110",
						 "000100011111110011000010",
						 "000100011111110110100110",
						 "000100011111111010001010",
						 "000100011111111101101110",
						 "000100100000000001010010",
						 "000100100000000100110110",
						 "000100100000001000011010",
						 "000100100000001011111110",
						 "000100100000001111100010",
						 "000100100000010011000110",
						 "000100100000010110101010",
						 "000100100000011010001110",
						 "000100100000011101110010",
						 "000100100000100001010110",
						 "000100100000100100111010",
						 "000100100010010010011100",
						 "000100100010010110000000",
						 "000100100010011001100100",
						 "000100100010011101001000",
						 "000100100010100000101100",
						 "000100100010100100010000",
						 "000100100010100111110100",
						 "000100100010101011011000",
						 "000100100010101110111100",
						 "000100100010110010100000",
						 "000100100010110110000100",
						 "000100100010111001101000",
						 "000100100010111101001100",
						 "000100100011000000110000",
						 "000100100011000100010100",
						 "000100100011000111111000",
						 "000100100010010010011100",
						 "000100100010010110000000",
						 "000100100010011001100100",
						 "000100100010011101001000",
						 "000100100010100000101100",
						 "000100100010100100010000",
						 "000100100010100111110100",
						 "000100100010101011011000",
						 "000100100010101110111100",
						 "000100100010110010100000",
						 "000100100010110110000100",
						 "000100100010111001101000",
						 "000100100010111101001100",
						 "000100100011000000110000",
						 "000100100011000100010100",
						 "000100100011000111111000",
						 "000100100010010010011100",
						 "000100100010010110000000",
						 "000100100010011001100100",
						 "000100100010011101001000",
						 "000100100010100000101100",
						 "000100100010100100010000",
						 "000100100010100111110100",
						 "000100100010101011011000",
						 "000100100010101110111100",
						 "000100100010110010100000",
						 "000100100010110110000100",
						 "000100100010111001101000",
						 "000100100010111101001100",
						 "000100100011000000110000",
						 "000100100011000100010100",
						 "000100100011000111111000",
						 "000100100100110101011010",
						 "000100100100111000111110",
						 "000100100100111100100010",
						 "000100100101000000000110",
						 "000100100101000011101010",
						 "000100100101000111001110",
						 "000100100101001010110010",
						 "000100100101001110010110",
						 "000100100101010001111010",
						 "000100100101010101011110",
						 "000100100101011001000010",
						 "000100100101011100100110",
						 "000100100101100000001010",
						 "000100100101100011101110",
						 "000100100101100111010010",
						 "000100100101101010110110",
						 "000100100100110101011010",
						 "000100100100111000111110",
						 "000100100100111100100010",
						 "000100100101000000000110",
						 "000100100101000011101010",
						 "000100100101000111001110",
						 "000100100101001010110010",
						 "000100100101001110010110",
						 "000100100101010001111010",
						 "000100100101010101011110",
						 "000100100101011001000010",
						 "000100100101011100100110",
						 "000100100101100000001010",
						 "000100100101100011101110",
						 "000100100101100111010010",
						 "000100100101101010110110",
						 "000100100100110101011010",
						 "000100100100111000111101",
						 "000100100100111100100000",
						 "000100100101000000000011",
						 "000100100101000011100110",
						 "000100100101000111001001",
						 "000100100101001010101100",
						 "000100100101001110001111",
						 "000100100101010001110010",
						 "000100100101010101010101",
						 "000100100101011000111000",
						 "000100100101011100011011",
						 "000100100101011111111110",
						 "000100100101100011100001",
						 "000100100101100111000100",
						 "000100100101101010100111",
						 "000100100111011000011000",
						 "000100100111011011111011",
						 "000100100111011111011110",
						 "000100100111100011000001",
						 "000100100111100110100100",
						 "000100100111101010000111",
						 "000100100111101101101010",
						 "000100100111110001001101",
						 "000100100111110100110000",
						 "000100100111111000010011",
						 "000100100111111011110110",
						 "000100100111111111011001",
						 "000100101000000010111100",
						 "000100101000000110011111",
						 "000100101000001010000010",
						 "000100101000001101100101",
						 "000100100111011000011000",
						 "000100100111011011111011",
						 "000100100111011111011110",
						 "000100100111100011000001",
						 "000100100111100110100100",
						 "000100100111101010000111",
						 "000100100111101101101010",
						 "000100100111110001001101",
						 "000100100111110100110000",
						 "000100100111111000010011",
						 "000100100111111011110110",
						 "000100100111111111011001",
						 "000100101000000010111100",
						 "000100101000000110011111",
						 "000100101000001010000010",
						 "000100101000001101100101",
						 "000100100111011000011000",
						 "000100100111011011111011",
						 "000100100111011111011110",
						 "000100100111100011000001",
						 "000100100111100110100100",
						 "000100100111101010000111",
						 "000100100111101101101010",
						 "000100100111110001001101",
						 "000100100111110100110000",
						 "000100100111111000010011",
						 "000100100111111011110110",
						 "000100100111111111011001",
						 "000100101000000010111100",
						 "000100101000000110011111",
						 "000100101000001010000010",
						 "000100101000001101100101",
						 "000100101001111011010110",
						 "000100101001111110111001",
						 "000100101010000010011100",
						 "000100101010000101111111",
						 "000100101010001001100010",
						 "000100101010001101000101",
						 "000100101010010000101000",
						 "000100101010010100001011",
						 "000100101010010111101110",
						 "000100101010011011010001",
						 "000100101010011110110100",
						 "000100101010100010010111",
						 "000100101010100101111010",
						 "000100101010101001011101",
						 "000100101010101101000000",
						 "000100101010110000100011",
						 "000100101001111011010110",
						 "000100101001111110111000",
						 "000100101010000010011010",
						 "000100101010000101111100",
						 "000100101010001001011110",
						 "000100101010001101000000",
						 "000100101010010000100010",
						 "000100101010010100000100",
						 "000100101010010111100110",
						 "000100101010011011001000",
						 "000100101010011110101010",
						 "000100101010100010001100",
						 "000100101010100101101110",
						 "000100101010101001010000",
						 "000100101010101100110010",
						 "000100101010110000010100",
						 "000100101001111011010110",
						 "000100101001111110111000",
						 "000100101010000010011010",
						 "000100101010000101111100",
						 "000100101010001001011110",
						 "000100101010001101000000",
						 "000100101010010000100010",
						 "000100101010010100000100",
						 "000100101010010111100110",
						 "000100101010011011001000",
						 "000100101010011110101010",
						 "000100101010100010001100",
						 "000100101010100101101110",
						 "000100101010101001010000",
						 "000100101010101100110010",
						 "000100101010110000010100",
						 "000100101100011110010100",
						 "000100101100100001110110",
						 "000100101100100101011000",
						 "000100101100101000111010",
						 "000100101100101100011100",
						 "000100101100101111111110",
						 "000100101100110011100000",
						 "000100101100110111000010",
						 "000100101100111010100100",
						 "000100101100111110000110",
						 "000100101101000001101000",
						 "000100101101000101001010",
						 "000100101101001000101100",
						 "000100101101001100001110",
						 "000100101101001111110000",
						 "000100101101010011010010",
						 "000100101100011110010100",
						 "000100101100100001110110",
						 "000100101100100101011000",
						 "000100101100101000111010",
						 "000100101100101100011100",
						 "000100101100101111111110",
						 "000100101100110011100000",
						 "000100101100110111000010",
						 "000100101100111010100100",
						 "000100101100111110000110",
						 "000100101101000001101000",
						 "000100101101000101001010",
						 "000100101101001000101100",
						 "000100101101001100001110",
						 "000100101101001111110000",
						 "000100101101010011010010",
						 "000100101100011110010100",
						 "000100101100100001110110",
						 "000100101100100101011000",
						 "000100101100101000111010",
						 "000100101100101100011100",
						 "000100101100101111111110",
						 "000100101100110011100000",
						 "000100101100110111000010",
						 "000100101100111010100100",
						 "000100101100111110000110",
						 "000100101101000001101000",
						 "000100101101000101001010",
						 "000100101101001000101100",
						 "000100101101001100001110",
						 "000100101101001111110000",
						 "000100101101010011010010",
						 "000100101111000001010010",
						 "000100101111000100110100",
						 "000100101111001000010110",
						 "000100101111001011111000",
						 "000100101111001111011010",
						 "000100101111010010111100",
						 "000100101111010110011110",
						 "000100101111011010000000",
						 "000100101111011101100010",
						 "000100101111100001000100",
						 "000100101111100100100110",
						 "000100101111101000001000",
						 "000100101111101011101010",
						 "000100101111101111001100",
						 "000100101111110010101110",
						 "000100101111110110010000",
						 "000100101111000001010010",
						 "000100101111000100110011",
						 "000100101111001000010100",
						 "000100101111001011110101",
						 "000100101111001111010110",
						 "000100101111010010110111",
						 "000100101111010110011000",
						 "000100101111011001111001",
						 "000100101111011101011010",
						 "000100101111100000111011",
						 "000100101111100100011100",
						 "000100101111100111111101",
						 "000100101111101011011110",
						 "000100101111101110111111",
						 "000100101111110010100000",
						 "000100101111110110000001",
						 "000100110001100100010000",
						 "000100110001100111110001",
						 "000100110001101011010010",
						 "000100110001101110110011",
						 "000100110001110010010100",
						 "000100110001110101110101",
						 "000100110001111001010110",
						 "000100110001111100110111",
						 "000100110010000000011000",
						 "000100110010000011111001",
						 "000100110010000111011010",
						 "000100110010001010111011",
						 "000100110010001110011100",
						 "000100110010010001111101",
						 "000100110010010101011110",
						 "000100110010011000111111",
						 "000100110001100100010000",
						 "000100110001100111110001",
						 "000100110001101011010010",
						 "000100110001101110110011",
						 "000100110001110010010100",
						 "000100110001110101110101",
						 "000100110001111001010110",
						 "000100110001111100110111",
						 "000100110010000000011000",
						 "000100110010000011111001",
						 "000100110010000111011010",
						 "000100110010001010111011",
						 "000100110010001110011100",
						 "000100110010010001111101",
						 "000100110010010101011110",
						 "000100110010011000111111",
						 "000100110001100100010000",
						 "000100110001100111110001",
						 "000100110001101011010010",
						 "000100110001101110110011",
						 "000100110001110010010100",
						 "000100110001110101110101",
						 "000100110001111001010110",
						 "000100110001111100110111",
						 "000100110010000000011000",
						 "000100110010000011111001",
						 "000100110010000111011010",
						 "000100110010001010111011",
						 "000100110010001110011100",
						 "000100110010010001111101",
						 "000100110010010101011110",
						 "000100110010011000111111",
						 "000100110100000111001110",
						 "000100110100001010101111",
						 "000100110100001110010000",
						 "000100110100010001110001",
						 "000100110100010101010010",
						 "000100110100011000110011",
						 "000100110100011100010100",
						 "000100110100011111110101",
						 "000100110100100011010110",
						 "000100110100100110110111",
						 "000100110100101010011000",
						 "000100110100101101111001",
						 "000100110100110001011010",
						 "000100110100110100111011",
						 "000100110100111000011100",
						 "000100110100111011111101",
						 "000100110100000111001110",
						 "000100110100001010101110",
						 "000100110100001110001110",
						 "000100110100010001101110",
						 "000100110100010101001110",
						 "000100110100011000101110",
						 "000100110100011100001110",
						 "000100110100011111101110",
						 "000100110100100011001110",
						 "000100110100100110101110",
						 "000100110100101010001110",
						 "000100110100101101101110",
						 "000100110100110001001110",
						 "000100110100110100101110",
						 "000100110100111000001110",
						 "000100110100111011101110",
						 "000100110100000111001110",
						 "000100110100001010101110",
						 "000100110100001110001110",
						 "000100110100010001101110",
						 "000100110100010101001110",
						 "000100110100011000101110",
						 "000100110100011100001110",
						 "000100110100011111101110",
						 "000100110100100011001110",
						 "000100110100100110101110",
						 "000100110100101010001110",
						 "000100110100101101101110",
						 "000100110100110001001110",
						 "000100110100110100101110",
						 "000100110100111000001110",
						 "000100110100111011101110",
						 "000100110110101010001100",
						 "000100110110101101101100",
						 "000100110110110001001100",
						 "000100110110110100101100",
						 "000100110110111000001100",
						 "000100110110111011101100",
						 "000100110110111111001100",
						 "000100110111000010101100",
						 "000100110111000110001100",
						 "000100110111001001101100",
						 "000100110111001101001100",
						 "000100110111010000101100",
						 "000100110111010100001100",
						 "000100110111010111101100",
						 "000100110111011011001100",
						 "000100110111011110101100",
						 "000100110110101010001100",
						 "000100110110101101101100",
						 "000100110110110001001100",
						 "000100110110110100101100",
						 "000100110110111000001100",
						 "000100110110111011101100",
						 "000100110110111111001100",
						 "000100110111000010101100",
						 "000100110111000110001100",
						 "000100110111001001101100",
						 "000100110111001101001100",
						 "000100110111010000101100",
						 "000100110111010100001100",
						 "000100110111010111101100",
						 "000100110111011011001100",
						 "000100110111011110101100",
						 "000100110110101010001100",
						 "000100110110101101101100",
						 "000100110110110001001100",
						 "000100110110110100101100",
						 "000100110110111000001100",
						 "000100110110111011101100",
						 "000100110110111111001100",
						 "000100110111000010101100",
						 "000100110111000110001100",
						 "000100110111001001101100",
						 "000100110111001101001100",
						 "000100110111010000101100",
						 "000100110111010100001100",
						 "000100110111010111101100",
						 "000100110111011011001100",
						 "000100110111011110101100",
						 "000100111001001101001010",
						 "000100111001010000101001",
						 "000100111001010100001000",
						 "000100111001010111100111",
						 "000100111001011011000110",
						 "000100111001011110100101",
						 "000100111001100010000100",
						 "000100111001100101100011",
						 "000100111001101001000010",
						 "000100111001101100100001",
						 "000100111001110000000000",
						 "000100111001110011011111",
						 "000100111001110110111110",
						 "000100111001111010011101",
						 "000100111001111101111100",
						 "000100111010000001011011",
						 "000100111001001101001010",
						 "000100111001010000101001",
						 "000100111001010100001000",
						 "000100111001010111100111",
						 "000100111001011011000110",
						 "000100111001011110100101",
						 "000100111001100010000100",
						 "000100111001100101100011",
						 "000100111001101001000010",
						 "000100111001101100100001",
						 "000100111001110000000000",
						 "000100111001110011011111",
						 "000100111001110110111110",
						 "000100111001111010011101",
						 "000100111001111101111100",
						 "000100111010000001011011",
						 "000100111001001101001010",
						 "000100111001010000101001",
						 "000100111001010100001000",
						 "000100111001010111100111",
						 "000100111001011011000110",
						 "000100111001011110100101",
						 "000100111001100010000100",
						 "000100111001100101100011",
						 "000100111001101001000010",
						 "000100111001101100100001",
						 "000100111001110000000000",
						 "000100111001110011011111",
						 "000100111001110110111110",
						 "000100111001111010011101",
						 "000100111001111101111100",
						 "000100111010000001011011",
						 "000100111011110000001000",
						 "000100111011110011100111",
						 "000100111011110111000110",
						 "000100111011111010100101",
						 "000100111011111110000100",
						 "000100111100000001100011",
						 "000100111100000101000010",
						 "000100111100001000100001",
						 "000100111100001100000000",
						 "000100111100001111011111",
						 "000100111100010010111110",
						 "000100111100010110011101",
						 "000100111100011001111100",
						 "000100111100011101011011",
						 "000100111100100000111010",
						 "000100111100100100011001",
						 "000100111011110000001000",
						 "000100111011110011100111",
						 "000100111011110111000110",
						 "000100111011111010100101",
						 "000100111011111110000100",
						 "000100111100000001100011",
						 "000100111100000101000010",
						 "000100111100001000100001",
						 "000100111100001100000000",
						 "000100111100001111011111",
						 "000100111100010010111110",
						 "000100111100010110011101",
						 "000100111100011001111100",
						 "000100111100011101011011",
						 "000100111100100000111010",
						 "000100111100100100011001",
						 "000100111011110000001000",
						 "000100111011110011100111",
						 "000100111011110111000110",
						 "000100111011111010100101",
						 "000100111011111110000100",
						 "000100111100000001100011",
						 "000100111100000101000010",
						 "000100111100001000100001",
						 "000100111100001100000000",
						 "000100111100001111011111",
						 "000100111100010010111110",
						 "000100111100010110011101",
						 "000100111100011001111100",
						 "000100111100011101011011",
						 "000100111100100000111010",
						 "000100111100100100011001",
						 "000100111110010011000110",
						 "000100111110010110100100",
						 "000100111110011010000010",
						 "000100111110011101100000",
						 "000100111110100000111110",
						 "000100111110100100011100",
						 "000100111110100111111010",
						 "000100111110101011011000",
						 "000100111110101110110110",
						 "000100111110110010010100",
						 "000100111110110101110010",
						 "000100111110111001010000",
						 "000100111110111100101110",
						 "000100111111000000001100",
						 "000100111111000011101010",
						 "000100111111000111001000",
						 "000100111110010011000110",
						 "000100111110010110100100",
						 "000100111110011010000010",
						 "000100111110011101100000",
						 "000100111110100000111110",
						 "000100111110100100011100",
						 "000100111110100111111010",
						 "000100111110101011011000",
						 "000100111110101110110110",
						 "000100111110110010010100",
						 "000100111110110101110010",
						 "000100111110111001010000",
						 "000100111110111100101110",
						 "000100111111000000001100",
						 "000100111111000011101010",
						 "000100111111000111001000",
						 "000100111110010011000110",
						 "000100111110010110100100",
						 "000100111110011010000010",
						 "000100111110011101100000",
						 "000100111110100000111110",
						 "000100111110100100011100",
						 "000100111110100111111010",
						 "000100111110101011011000",
						 "000100111110101110110110",
						 "000100111110110010010100",
						 "000100111110110101110010",
						 "000100111110111001010000",
						 "000100111110111100101110",
						 "000100111111000000001100",
						 "000100111111000011101010",
						 "000100111111000111001000",
						 "000101000000110110000100",
						 "000101000000111001100010",
						 "000101000000111101000000",
						 "000101000001000000011110",
						 "000101000001000011111100",
						 "000101000001000111011010",
						 "000101000001001010111000",
						 "000101000001001110010110",
						 "000101000001010001110100",
						 "000101000001010101010010",
						 "000101000001011000110000",
						 "000101000001011100001110",
						 "000101000001011111101100",
						 "000101000001100011001010",
						 "000101000001100110101000",
						 "000101000001101010000110",
						 "000101000000110110000100",
						 "000101000000111001100010",
						 "000101000000111101000000",
						 "000101000001000000011110",
						 "000101000001000011111100",
						 "000101000001000111011010",
						 "000101000001001010111000",
						 "000101000001001110010110",
						 "000101000001010001110100",
						 "000101000001010101010010",
						 "000101000001011000110000",
						 "000101000001011100001110",
						 "000101000001011111101100",
						 "000101000001100011001010",
						 "000101000001100110101000",
						 "000101000001101010000110",
						 "000101000000110110000100",
						 "000101000000111001100001",
						 "000101000000111100111110",
						 "000101000001000000011011",
						 "000101000001000011111000",
						 "000101000001000111010101",
						 "000101000001001010110010",
						 "000101000001001110001111",
						 "000101000001010001101100",
						 "000101000001010101001001",
						 "000101000001011000100110",
						 "000101000001011100000011",
						 "000101000001011111100000",
						 "000101000001100010111101",
						 "000101000001100110011010",
						 "000101000001101001110111",
						 "000101000011011001000010",
						 "000101000011011100011111",
						 "000101000011011111111100",
						 "000101000011100011011001",
						 "000101000011100110110110",
						 "000101000011101010010011",
						 "000101000011101101110000",
						 "000101000011110001001101",
						 "000101000011110100101010",
						 "000101000011111000000111",
						 "000101000011111011100100",
						 "000101000011111111000001",
						 "000101000100000010011110",
						 "000101000100000101111011",
						 "000101000100001001011000",
						 "000101000100001100110101",
						 "000101000011011001000010",
						 "000101000011011100011111",
						 "000101000011011111111100",
						 "000101000011100011011001",
						 "000101000011100110110110",
						 "000101000011101010010011",
						 "000101000011101101110000",
						 "000101000011110001001101",
						 "000101000011110100101010",
						 "000101000011111000000111",
						 "000101000011111011100100",
						 "000101000011111111000001",
						 "000101000100000010011110",
						 "000101000100000101111011",
						 "000101000100001001011000",
						 "000101000100001100110101",
						 "000101000011011001000010",
						 "000101000011011100011111",
						 "000101000011011111111100",
						 "000101000011100011011001",
						 "000101000011100110110110",
						 "000101000011101010010011",
						 "000101000011101101110000",
						 "000101000011110001001101",
						 "000101000011110100101010",
						 "000101000011111000000111",
						 "000101000011111011100100",
						 "000101000011111111000001",
						 "000101000100000010011110",
						 "000101000100000101111011",
						 "000101000100001001011000",
						 "000101000100001100110101",
						 "000101000101111100000000",
						 "000101000101111111011101",
						 "000101000110000010111010",
						 "000101000110000110010111",
						 "000101000110001001110100",
						 "000101000110001101010001",
						 "000101000110010000101110",
						 "000101000110010100001011",
						 "000101000110010111101000",
						 "000101000110011011000101",
						 "000101000110011110100010",
						 "000101000110100001111111",
						 "000101000110100101011100",
						 "000101000110101000111001",
						 "000101000110101100010110",
						 "000101000110101111110011",
						 "000101000101111100000000",
						 "000101000101111111011100",
						 "000101000110000010111000",
						 "000101000110000110010100",
						 "000101000110001001110000",
						 "000101000110001101001100",
						 "000101000110010000101000",
						 "000101000110010100000100",
						 "000101000110010111100000",
						 "000101000110011010111100",
						 "000101000110011110011000",
						 "000101000110100001110100",
						 "000101000110100101010000",
						 "000101000110101000101100",
						 "000101000110101100001000",
						 "000101000110101111100100",
						 "000101000101111100000000",
						 "000101000101111111011100",
						 "000101000110000010111000",
						 "000101000110000110010100",
						 "000101000110001001110000",
						 "000101000110001101001100",
						 "000101000110010000101000",
						 "000101000110010100000100",
						 "000101000110010111100000",
						 "000101000110011010111100",
						 "000101000110011110011000",
						 "000101000110100001110100",
						 "000101000110100101010000",
						 "000101000110101000101100",
						 "000101000110101100001000",
						 "000101000110101111100100",
						 "000101001000011110111110",
						 "000101001000100010011010",
						 "000101001000100101110110",
						 "000101001000101001010010",
						 "000101001000101100101110",
						 "000101001000110000001010",
						 "000101001000110011100110",
						 "000101001000110111000010",
						 "000101001000111010011110",
						 "000101001000111101111010",
						 "000101001001000001010110",
						 "000101001001000100110010",
						 "000101001001001000001110",
						 "000101001001001011101010",
						 "000101001001001111000110",
						 "000101001001010010100010",
						 "000101001000011110111110",
						 "000101001000100010011010",
						 "000101001000100101110110",
						 "000101001000101001010010",
						 "000101001000101100101110",
						 "000101001000110000001010",
						 "000101001000110011100110",
						 "000101001000110111000010",
						 "000101001000111010011110",
						 "000101001000111101111010",
						 "000101001001000001010110",
						 "000101001001000100110010",
						 "000101001001001000001110",
						 "000101001001001011101010",
						 "000101001001001111000110",
						 "000101001001010010100010",
						 "000101001000011110111110",
						 "000101001000100010011010",
						 "000101001000100101110110",
						 "000101001000101001010010",
						 "000101001000101100101110",
						 "000101001000110000001010",
						 "000101001000110011100110",
						 "000101001000110111000010",
						 "000101001000111010011110",
						 "000101001000111101111010",
						 "000101001001000001010110",
						 "000101001001000100110010",
						 "000101001001001000001110",
						 "000101001001001011101010",
						 "000101001001001111000110",
						 "000101001001010010100010",
						 "000101001011000001111100",
						 "000101001011000101010111",
						 "000101001011001000110010",
						 "000101001011001100001101",
						 "000101001011001111101000",
						 "000101001011010011000011",
						 "000101001011010110011110",
						 "000101001011011001111001",
						 "000101001011011101010100",
						 "000101001011100000101111",
						 "000101001011100100001010",
						 "000101001011100111100101",
						 "000101001011101011000000",
						 "000101001011101110011011",
						 "000101001011110001110110",
						 "000101001011110101010001",
						 "000101001011000001111100",
						 "000101001011000101010111",
						 "000101001011001000110010",
						 "000101001011001100001101",
						 "000101001011001111101000",
						 "000101001011010011000011",
						 "000101001011010110011110",
						 "000101001011011001111001",
						 "000101001011011101010100",
						 "000101001011100000101111",
						 "000101001011100100001010",
						 "000101001011100111100101",
						 "000101001011101011000000",
						 "000101001011101110011011",
						 "000101001011110001110110",
						 "000101001011110101010001",
						 "000101001011000001111100",
						 "000101001011000101010111",
						 "000101001011001000110010",
						 "000101001011001100001101",
						 "000101001011001111101000",
						 "000101001011010011000011",
						 "000101001011010110011110",
						 "000101001011011001111001",
						 "000101001011011101010100",
						 "000101001011100000101111",
						 "000101001011100100001010",
						 "000101001011100111100101",
						 "000101001011101011000000",
						 "000101001011101110011011",
						 "000101001011110001110110",
						 "000101001011110101010001",
						 "000101001101100100111010",
						 "000101001101101000010101",
						 "000101001101101011110000",
						 "000101001101101111001011",
						 "000101001101110010100110",
						 "000101001101110110000001",
						 "000101001101111001011100",
						 "000101001101111100110111",
						 "000101001110000000010010",
						 "000101001110000011101101",
						 "000101001110000111001000",
						 "000101001110001010100011",
						 "000101001110001101111110",
						 "000101001110010001011001",
						 "000101001110010100110100",
						 "000101001110011000001111",
						 "000101001101100100111010",
						 "000101001101101000010101",
						 "000101001101101011110000",
						 "000101001101101111001011",
						 "000101001101110010100110",
						 "000101001101110110000001",
						 "000101001101111001011100",
						 "000101001101111100110111",
						 "000101001110000000010010",
						 "000101001110000011101101",
						 "000101001110000111001000",
						 "000101001110001010100011",
						 "000101001110001101111110",
						 "000101001110010001011001",
						 "000101001110010100110100",
						 "000101001110011000001111",
						 "000101001101100100111010",
						 "000101001101101000010100",
						 "000101001101101011101110",
						 "000101001101101111001000",
						 "000101001101110010100010",
						 "000101001101110101111100",
						 "000101001101111001010110",
						 "000101001101111100110000",
						 "000101001110000000001010",
						 "000101001110000011100100",
						 "000101001110000110111110",
						 "000101001110001010011000",
						 "000101001110001101110010",
						 "000101001110010001001100",
						 "000101001110010100100110",
						 "000101001110011000000000",
						 "000101010000000111111000",
						 "000101010000001011010010",
						 "000101010000001110101100",
						 "000101010000010010000110",
						 "000101010000010101100000",
						 "000101010000011000111010",
						 "000101010000011100010100",
						 "000101010000011111101110",
						 "000101010000100011001000",
						 "000101010000100110100010",
						 "000101010000101001111100",
						 "000101010000101101010110",
						 "000101010000110000110000",
						 "000101010000110100001010",
						 "000101010000110111100100",
						 "000101010000111010111110",
						 "000101010000000111111000",
						 "000101010000001011010010",
						 "000101010000001110101100",
						 "000101010000010010000110",
						 "000101010000010101100000",
						 "000101010000011000111010",
						 "000101010000011100010100",
						 "000101010000011111101110",
						 "000101010000100011001000",
						 "000101010000100110100010",
						 "000101010000101001111100",
						 "000101010000101101010110",
						 "000101010000110000110000",
						 "000101010000110100001010",
						 "000101010000110111100100",
						 "000101010000111010111110",
						 "000101010000000111111000",
						 "000101010000001011010010",
						 "000101010000001110101100",
						 "000101010000010010000110",
						 "000101010000010101100000",
						 "000101010000011000111010",
						 "000101010000011100010100",
						 "000101010000011111101110",
						 "000101010000100011001000",
						 "000101010000100110100010",
						 "000101010000101001111100",
						 "000101010000101101010110",
						 "000101010000110000110000",
						 "000101010000110100001010",
						 "000101010000110111100100",
						 "000101010000111010111110",
						 "000101010010101010110110",
						 "000101010010101110010000",
						 "000101010010110001101010",
						 "000101010010110101000100",
						 "000101010010111000011110",
						 "000101010010111011111000",
						 "000101010010111111010010",
						 "000101010011000010101100",
						 "000101010011000110000110",
						 "000101010011001001100000",
						 "000101010011001100111010",
						 "000101010011010000010100",
						 "000101010011010011101110",
						 "000101010011010111001000",
						 "000101010011011010100010",
						 "000101010011011101111100",
						 "000101010010101010110110",
						 "000101010010101110001111",
						 "000101010010110001101000",
						 "000101010010110101000001",
						 "000101010010111000011010",
						 "000101010010111011110011",
						 "000101010010111111001100",
						 "000101010011000010100101",
						 "000101010011000101111110",
						 "000101010011001001010111",
						 "000101010011001100110000",
						 "000101010011010000001001",
						 "000101010011010011100010",
						 "000101010011010110111011",
						 "000101010011011010010100",
						 "000101010011011101101101",
						 "000101010010101010110110",
						 "000101010010101110001111",
						 "000101010010110001101000",
						 "000101010010110101000001",
						 "000101010010111000011010",
						 "000101010010111011110011",
						 "000101010010111111001100",
						 "000101010011000010100101",
						 "000101010011000101111110",
						 "000101010011001001010111",
						 "000101010011001100110000",
						 "000101010011010000001001",
						 "000101010011010011100010",
						 "000101010011010110111011",
						 "000101010011011010010100",
						 "000101010011011101101101",
						 "000101010101001101110100",
						 "000101010101010001001101",
						 "000101010101010100100110",
						 "000101010101010111111111",
						 "000101010101011011011000",
						 "000101010101011110110001",
						 "000101010101100010001010",
						 "000101010101100101100011",
						 "000101010101101000111100",
						 "000101010101101100010101",
						 "000101010101101111101110",
						 "000101010101110011000111",
						 "000101010101110110100000",
						 "000101010101111001111001",
						 "000101010101111101010010",
						 "000101010110000000101011",
						 "000101010101001101110100",
						 "000101010101010001001101",
						 "000101010101010100100110",
						 "000101010101010111111111",
						 "000101010101011011011000",
						 "000101010101011110110001",
						 "000101010101100010001010",
						 "000101010101100101100011",
						 "000101010101101000111100",
						 "000101010101101100010101",
						 "000101010101101111101110",
						 "000101010101110011000111",
						 "000101010101110110100000",
						 "000101010101111001111001",
						 "000101010101111101010010",
						 "000101010110000000101011",
						 "000101010101001101110100",
						 "000101010101010001001101",
						 "000101010101010100100110",
						 "000101010101010111111111",
						 "000101010101011011011000",
						 "000101010101011110110001",
						 "000101010101100010001010",
						 "000101010101100101100011",
						 "000101010101101000111100",
						 "000101010101101100010101",
						 "000101010101101111101110",
						 "000101010101110011000111",
						 "000101010101110110100000",
						 "000101010101111001111001",
						 "000101010101111101010010",
						 "000101010110000000101011",
						 "000101010111110000110010",
						 "000101010111110100001010",
						 "000101010111110111100010",
						 "000101010111111010111010",
						 "000101010111111110010010",
						 "000101011000000001101010",
						 "000101011000000101000010",
						 "000101011000001000011010",
						 "000101011000001011110010",
						 "000101011000001111001010",
						 "000101011000010010100010",
						 "000101011000010101111010",
						 "000101011000011001010010",
						 "000101011000011100101010",
						 "000101011000100000000010",
						 "000101011000100011011010",
						 "000101010111110000110010",
						 "000101010111110100001010",
						 "000101010111110111100010",
						 "000101010111111010111010",
						 "000101010111111110010010",
						 "000101011000000001101010",
						 "000101011000000101000010",
						 "000101011000001000011010",
						 "000101011000001011110010",
						 "000101011000001111001010",
						 "000101011000010010100010",
						 "000101011000010101111010",
						 "000101011000011001010010",
						 "000101011000011100101010",
						 "000101011000100000000010",
						 "000101011000100011011010",
						 "000101010111110000110010",
						 "000101010111110100001010",
						 "000101010111110111100010",
						 "000101010111111010111010",
						 "000101010111111110010010",
						 "000101011000000001101010",
						 "000101011000000101000010",
						 "000101011000001000011010",
						 "000101011000001011110010",
						 "000101011000001111001010",
						 "000101011000010010100010",
						 "000101011000010101111010",
						 "000101011000011001010010",
						 "000101011000011100101010",
						 "000101011000100000000010",
						 "000101011000100011011010",
						 "000101011010010011110000",
						 "000101011010010111001000",
						 "000101011010011010100000",
						 "000101011010011101111000",
						 "000101011010100001010000",
						 "000101011010100100101000",
						 "000101011010101000000000",
						 "000101011010101011011000",
						 "000101011010101110110000",
						 "000101011010110010001000",
						 "000101011010110101100000",
						 "000101011010111000111000",
						 "000101011010111100010000",
						 "000101011010111111101000",
						 "000101011011000011000000",
						 "000101011011000110011000",
						 "000101011010010011110000",
						 "000101011010010111001000",
						 "000101011010011010100000",
						 "000101011010011101111000",
						 "000101011010100001010000",
						 "000101011010100100101000",
						 "000101011010101000000000",
						 "000101011010101011011000",
						 "000101011010101110110000",
						 "000101011010110010001000",
						 "000101011010110101100000",
						 "000101011010111000111000",
						 "000101011010111100010000",
						 "000101011010111111101000",
						 "000101011011000011000000",
						 "000101011011000110011000",
						 "000101011010010011110000",
						 "000101011010010111000111",
						 "000101011010011010011110",
						 "000101011010011101110101",
						 "000101011010100001001100",
						 "000101011010100100100011",
						 "000101011010100111111010",
						 "000101011010101011010001",
						 "000101011010101110101000",
						 "000101011010110001111111",
						 "000101011010110101010110",
						 "000101011010111000101101",
						 "000101011010111100000100",
						 "000101011010111111011011",
						 "000101011011000010110010",
						 "000101011011000110001001",
						 "000101011100110110101110",
						 "000101011100111010000101",
						 "000101011100111101011100",
						 "000101011101000000110011",
						 "000101011101000100001010",
						 "000101011101000111100001",
						 "000101011101001010111000",
						 "000101011101001110001111",
						 "000101011101010001100110",
						 "000101011101010100111101",
						 "000101011101011000010100",
						 "000101011101011011101011",
						 "000101011101011111000010",
						 "000101011101100010011001",
						 "000101011101100101110000",
						 "000101011101101001000111",
						 "000101011100110110101110",
						 "000101011100111010000101",
						 "000101011100111101011100",
						 "000101011101000000110011",
						 "000101011101000100001010",
						 "000101011101000111100001",
						 "000101011101001010111000",
						 "000101011101001110001111",
						 "000101011101010001100110",
						 "000101011101010100111101",
						 "000101011101011000010100",
						 "000101011101011011101011",
						 "000101011101011111000010",
						 "000101011101100010011001",
						 "000101011101100101110000",
						 "000101011101101001000111",
						 "000101011100110110101110",
						 "000101011100111010000101",
						 "000101011100111101011100",
						 "000101011101000000110011",
						 "000101011101000100001010",
						 "000101011101000111100001",
						 "000101011101001010111000",
						 "000101011101001110001111",
						 "000101011101010001100110",
						 "000101011101010100111101",
						 "000101011101011000010100",
						 "000101011101011011101011",
						 "000101011101011111000010",
						 "000101011101100010011001",
						 "000101011101100101110000",
						 "000101011101101001000111",
						 "000101011111011001101100",
						 "000101011111011101000010",
						 "000101011111100000011000",
						 "000101011111100011101110",
						 "000101011111100111000100",
						 "000101011111101010011010",
						 "000101011111101101110000",
						 "000101011111110001000110",
						 "000101011111110100011100",
						 "000101011111110111110010",
						 "000101011111111011001000",
						 "000101011111111110011110",
						 "000101100000000001110100",
						 "000101100000000101001010",
						 "000101100000001000100000",
						 "000101100000001011110110",
						 "000101011111011001101100",
						 "000101011111011101000010",
						 "000101011111100000011000",
						 "000101011111100011101110",
						 "000101011111100111000100",
						 "000101011111101010011010",
						 "000101011111101101110000",
						 "000101011111110001000110",
						 "000101011111110100011100",
						 "000101011111110111110010",
						 "000101011111111011001000",
						 "000101011111111110011110",
						 "000101100000000001110100",
						 "000101100000000101001010",
						 "000101100000001000100000",
						 "000101100000001011110110",
						 "000101011111011001101100",
						 "000101011111011101000010",
						 "000101011111100000011000",
						 "000101011111100011101110",
						 "000101011111100111000100",
						 "000101011111101010011010",
						 "000101011111101101110000",
						 "000101011111110001000110",
						 "000101011111110100011100",
						 "000101011111110111110010",
						 "000101011111111011001000",
						 "000101011111111110011110",
						 "000101100000000001110100",
						 "000101100000000101001010",
						 "000101100000001000100000",
						 "000101100000001011110110",
						 "000101100001111100101010",
						 "000101100010000000000000",
						 "000101100010000011010110",
						 "000101100010000110101100",
						 "000101100010001010000010",
						 "000101100010001101011000",
						 "000101100010010000101110",
						 "000101100010010100000100",
						 "000101100010010111011010",
						 "000101100010011010110000",
						 "000101100010011110000110",
						 "000101100010100001011100",
						 "000101100010100100110010",
						 "000101100010101000001000",
						 "000101100010101011011110",
						 "000101100010101110110100",
						 "000101100001111100101010",
						 "000101100010000000000000",
						 "000101100010000011010110",
						 "000101100010000110101100",
						 "000101100010001010000010",
						 "000101100010001101011000",
						 "000101100010010000101110",
						 "000101100010010100000100",
						 "000101100010010111011010",
						 "000101100010011010110000",
						 "000101100010011110000110",
						 "000101100010100001011100",
						 "000101100010100100110010",
						 "000101100010101000001000",
						 "000101100010101011011110",
						 "000101100010101110110100",
						 "000101100001111100101010",
						 "000101100001111111111111",
						 "000101100010000011010100",
						 "000101100010000110101001",
						 "000101100010001001111110",
						 "000101100010001101010011",
						 "000101100010010000101000",
						 "000101100010010011111101",
						 "000101100010010111010010",
						 "000101100010011010100111",
						 "000101100010011101111100",
						 "000101100010100001010001",
						 "000101100010100100100110",
						 "000101100010100111111011",
						 "000101100010101011010000",
						 "000101100010101110100101",
						 "000101100100011111101000",
						 "000101100100100010111101",
						 "000101100100100110010010",
						 "000101100100101001100111",
						 "000101100100101100111100",
						 "000101100100110000010001",
						 "000101100100110011100110",
						 "000101100100110110111011",
						 "000101100100111010010000",
						 "000101100100111101100101",
						 "000101100101000000111010",
						 "000101100101000100001111",
						 "000101100101000111100100",
						 "000101100101001010111001",
						 "000101100101001110001110",
						 "000101100101010001100011",
						 "000101100100011111101000",
						 "000101100100100010111101",
						 "000101100100100110010010",
						 "000101100100101001100111",
						 "000101100100101100111100",
						 "000101100100110000010001",
						 "000101100100110011100110",
						 "000101100100110110111011",
						 "000101100100111010010000",
						 "000101100100111101100101",
						 "000101100101000000111010",
						 "000101100101000100001111",
						 "000101100101000111100100",
						 "000101100101001010111001",
						 "000101100101001110001110",
						 "000101100101010001100011",
						 "000101100100011111101000",
						 "000101100100100010111101",
						 "000101100100100110010010",
						 "000101100100101001100111",
						 "000101100100101100111100",
						 "000101100100110000010001",
						 "000101100100110011100110",
						 "000101100100110110111011",
						 "000101100100111010010000",
						 "000101100100111101100101",
						 "000101100101000000111010",
						 "000101100101000100001111",
						 "000101100101000111100100",
						 "000101100101001010111001",
						 "000101100101001110001110",
						 "000101100101010001100011",
						 "000101100111000010100110",
						 "000101100111000101111011",
						 "000101100111001001010000",
						 "000101100111001100100101",
						 "000101100111001111111010",
						 "000101100111010011001111",
						 "000101100111010110100100",
						 "000101100111011001111001",
						 "000101100111011101001110",
						 "000101100111100000100011",
						 "000101100111100011111000",
						 "000101100111100111001101",
						 "000101100111101010100010",
						 "000101100111101101110111",
						 "000101100111110001001100",
						 "000101100111110100100001",
						 "000101100111000010100110",
						 "000101100111000101111010",
						 "000101100111001001001110",
						 "000101100111001100100010",
						 "000101100111001111110110",
						 "000101100111010011001010",
						 "000101100111010110011110",
						 "000101100111011001110010",
						 "000101100111011101000110",
						 "000101100111100000011010",
						 "000101100111100011101110",
						 "000101100111100111000010",
						 "000101100111101010010110",
						 "000101100111101101101010",
						 "000101100111110000111110",
						 "000101100111110100010010",
						 "000101100111000010100110",
						 "000101100111000101111010",
						 "000101100111001001001110",
						 "000101100111001100100010",
						 "000101100111001111110110",
						 "000101100111010011001010",
						 "000101100111010110011110",
						 "000101100111011001110010",
						 "000101100111011101000110",
						 "000101100111100000011010",
						 "000101100111100011101110",
						 "000101100111100111000010",
						 "000101100111101010010110",
						 "000101100111101101101010",
						 "000101100111110000111110",
						 "000101100111110100010010",
						 "000101101001100101100100",
						 "000101101001101000111000",
						 "000101101001101100001100",
						 "000101101001101111100000",
						 "000101101001110010110100",
						 "000101101001110110001000",
						 "000101101001111001011100",
						 "000101101001111100110000",
						 "000101101010000000000100",
						 "000101101010000011011000",
						 "000101101010000110101100",
						 "000101101010001010000000",
						 "000101101010001101010100",
						 "000101101010010000101000",
						 "000101101010010011111100",
						 "000101101010010111010000",
						 "000101101001100101100100",
						 "000101101001101000111000",
						 "000101101001101100001100",
						 "000101101001101111100000",
						 "000101101001110010110100",
						 "000101101001110110001000",
						 "000101101001111001011100",
						 "000101101001111100110000",
						 "000101101010000000000100",
						 "000101101010000011011000",
						 "000101101010000110101100",
						 "000101101010001010000000",
						 "000101101010001101010100",
						 "000101101010010000101000",
						 "000101101010010011111100",
						 "000101101010010111010000",
						 "000101101001100101100100",
						 "000101101001101000110111",
						 "000101101001101100001010",
						 "000101101001101111011101",
						 "000101101001110010110000",
						 "000101101001110110000011",
						 "000101101001111001010110",
						 "000101101001111100101001",
						 "000101101001111111111100",
						 "000101101010000011001111",
						 "000101101010000110100010",
						 "000101101010001001110101",
						 "000101101010001101001000",
						 "000101101010010000011011",
						 "000101101010010011101110",
						 "000101101010010111000001",
						 "000101101100001000100010",
						 "000101101100001011110101",
						 "000101101100001111001000",
						 "000101101100010010011011",
						 "000101101100010101101110",
						 "000101101100011001000001",
						 "000101101100011100010100",
						 "000101101100011111100111",
						 "000101101100100010111010",
						 "000101101100100110001101",
						 "000101101100101001100000",
						 "000101101100101100110011",
						 "000101101100110000000110",
						 "000101101100110011011001",
						 "000101101100110110101100",
						 "000101101100111001111111",
						 "000101101100001000100010",
						 "000101101100001011110101",
						 "000101101100001111001000",
						 "000101101100010010011011",
						 "000101101100010101101110",
						 "000101101100011001000001",
						 "000101101100011100010100",
						 "000101101100011111100111",
						 "000101101100100010111010",
						 "000101101100100110001101",
						 "000101101100101001100000",
						 "000101101100101100110011",
						 "000101101100110000000110",
						 "000101101100110011011001",
						 "000101101100110110101100",
						 "000101101100111001111111",
						 "000101101100001000100010",
						 "000101101100001011110101",
						 "000101101100001111001000",
						 "000101101100010010011011",
						 "000101101100010101101110",
						 "000101101100011001000001",
						 "000101101100011100010100",
						 "000101101100011111100111",
						 "000101101100100010111010",
						 "000101101100100110001101",
						 "000101101100101001100000",
						 "000101101100101100110011",
						 "000101101100110000000110",
						 "000101101100110011011001",
						 "000101101100110110101100",
						 "000101101100111001111111",
						 "000101101110101011100000",
						 "000101101110101110110011",
						 "000101101110110010000110",
						 "000101101110110101011001",
						 "000101101110111000101100",
						 "000101101110111011111111",
						 "000101101110111111010010",
						 "000101101111000010100101",
						 "000101101111000101111000",
						 "000101101111001001001011",
						 "000101101111001100011110",
						 "000101101111001111110001",
						 "000101101111010011000100",
						 "000101101111010110010111",
						 "000101101111011001101010",
						 "000101101111011100111101",
						 "000101101110101011100000",
						 "000101101110101110110010",
						 "000101101110110010000100",
						 "000101101110110101010110",
						 "000101101110111000101000",
						 "000101101110111011111010",
						 "000101101110111111001100",
						 "000101101111000010011110",
						 "000101101111000101110000",
						 "000101101111001001000010",
						 "000101101111001100010100",
						 "000101101111001111100110",
						 "000101101111010010111000",
						 "000101101111010110001010",
						 "000101101111011001011100",
						 "000101101111011100101110",
						 "000101101110101011100000",
						 "000101101110101110110010",
						 "000101101110110010000100",
						 "000101101110110101010110",
						 "000101101110111000101000",
						 "000101101110111011111010",
						 "000101101110111111001100",
						 "000101101111000010011110",
						 "000101101111000101110000",
						 "000101101111001001000010",
						 "000101101111001100010100",
						 "000101101111001111100110",
						 "000101101111010010111000",
						 "000101101111010110001010",
						 "000101101111011001011100",
						 "000101101111011100101110",
						 "000101110001001110011110",
						 "000101110001010001110000",
						 "000101110001010101000010",
						 "000101110001011000010100",
						 "000101110001011011100110",
						 "000101110001011110111000",
						 "000101110001100010001010",
						 "000101110001100101011100",
						 "000101110001101000101110",
						 "000101110001101100000000",
						 "000101110001101111010010",
						 "000101110001110010100100",
						 "000101110001110101110110",
						 "000101110001111001001000",
						 "000101110001111100011010",
						 "000101110001111111101100",
						 "000101110001001110011110",
						 "000101110001010001110000",
						 "000101110001010101000010",
						 "000101110001011000010100",
						 "000101110001011011100110",
						 "000101110001011110111000",
						 "000101110001100010001010",
						 "000101110001100101011100",
						 "000101110001101000101110",
						 "000101110001101100000000",
						 "000101110001101111010010",
						 "000101110001110010100100",
						 "000101110001110101110110",
						 "000101110001111001001000",
						 "000101110001111100011010",
						 "000101110001111111101100",
						 "000101110001001110011110",
						 "000101110001010001101111",
						 "000101110001010101000000",
						 "000101110001011000010001",
						 "000101110001011011100010",
						 "000101110001011110110011",
						 "000101110001100010000100",
						 "000101110001100101010101",
						 "000101110001101000100110",
						 "000101110001101011110111",
						 "000101110001101111001000",
						 "000101110001110010011001",
						 "000101110001110101101010",
						 "000101110001111000111011",
						 "000101110001111100001100",
						 "000101110001111111011101",
						 "000101110011110001011100",
						 "000101110011110100101101",
						 "000101110011110111111110",
						 "000101110011111011001111",
						 "000101110011111110100000",
						 "000101110100000001110001",
						 "000101110100000101000010",
						 "000101110100001000010011",
						 "000101110100001011100100",
						 "000101110100001110110101",
						 "000101110100010010000110",
						 "000101110100010101010111",
						 "000101110100011000101000",
						 "000101110100011011111001",
						 "000101110100011111001010",
						 "000101110100100010011011",
						 "000101110011110001011100",
						 "000101110011110100101101",
						 "000101110011110111111110",
						 "000101110011111011001111",
						 "000101110011111110100000",
						 "000101110100000001110001",
						 "000101110100000101000010",
						 "000101110100001000010011",
						 "000101110100001011100100",
						 "000101110100001110110101",
						 "000101110100010010000110",
						 "000101110100010101010111",
						 "000101110100011000101000",
						 "000101110100011011111001",
						 "000101110100011111001010",
						 "000101110100100010011011",
						 "000101110011110001011100",
						 "000101110011110100101101",
						 "000101110011110111111110",
						 "000101110011111011001111",
						 "000101110011111110100000",
						 "000101110100000001110001",
						 "000101110100000101000010",
						 "000101110100001000010011",
						 "000101110100001011100100",
						 "000101110100001110110101",
						 "000101110100010010000110",
						 "000101110100010101010111",
						 "000101110100011000101000",
						 "000101110100011011111001",
						 "000101110100011111001010",
						 "000101110100100010011011",
						 "000101110110010100011010",
						 "000101110110010111101011",
						 "000101110110011010111100",
						 "000101110110011110001101",
						 "000101110110100001011110",
						 "000101110110100100101111",
						 "000101110110101000000000",
						 "000101110110101011010001",
						 "000101110110101110100010",
						 "000101110110110001110011",
						 "000101110110110101000100",
						 "000101110110111000010101",
						 "000101110110111011100110",
						 "000101110110111110110111",
						 "000101110111000010001000",
						 "000101110111000101011001",
						 "000101110110010100011010",
						 "000101110110010111101010",
						 "000101110110011010111010",
						 "000101110110011110001010",
						 "000101110110100001011010",
						 "000101110110100100101010",
						 "000101110110100111111010",
						 "000101110110101011001010",
						 "000101110110101110011010",
						 "000101110110110001101010",
						 "000101110110110100111010",
						 "000101110110111000001010",
						 "000101110110111011011010",
						 "000101110110111110101010",
						 "000101110111000001111010",
						 "000101110111000101001010",
						 "000101110110010100011010",
						 "000101110110010111101010",
						 "000101110110011010111010",
						 "000101110110011110001010",
						 "000101110110100001011010",
						 "000101110110100100101010",
						 "000101110110100111111010",
						 "000101110110101011001010",
						 "000101110110101110011010",
						 "000101110110110001101010",
						 "000101110110110100111010",
						 "000101110110111000001010",
						 "000101110110111011011010",
						 "000101110110111110101010",
						 "000101110111000001111010",
						 "000101110111000101001010",
						 "000101110110010100011010",
						 "000101110110010111101010",
						 "000101110110011010111010",
						 "000101110110011110001010",
						 "000101110110100001011010",
						 "000101110110100100101010",
						 "000101110110100111111010",
						 "000101110110101011001010",
						 "000101110110101110011010",
						 "000101110110110001101010",
						 "000101110110110100111010",
						 "000101110110111000001010",
						 "000101110110111011011010",
						 "000101110110111110101010",
						 "000101110111000001111010",
						 "000101110111000101001010",
						 "000101111000110111011000",
						 "000101111000111010101000",
						 "000101111000111101111000",
						 "000101111001000001001000",
						 "000101111001000100011000",
						 "000101111001000111101000",
						 "000101111001001010111000",
						 "000101111001001110001000",
						 "000101111001010001011000",
						 "000101111001010100101000",
						 "000101111001010111111000",
						 "000101111001011011001000",
						 "000101111001011110011000",
						 "000101111001100001101000",
						 "000101111001100100111000",
						 "000101111001101000001000",
						 "000101111000110111011000",
						 "000101111000111010100111",
						 "000101111000111101110110",
						 "000101111001000001000101",
						 "000101111001000100010100",
						 "000101111001000111100011",
						 "000101111001001010110010",
						 "000101111001001110000001",
						 "000101111001010001010000",
						 "000101111001010100011111",
						 "000101111001010111101110",
						 "000101111001011010111101",
						 "000101111001011110001100",
						 "000101111001100001011011",
						 "000101111001100100101010",
						 "000101111001100111111001",
						 "000101111000110111011000",
						 "000101111000111010100111",
						 "000101111000111101110110",
						 "000101111001000001000101",
						 "000101111001000100010100",
						 "000101111001000111100011",
						 "000101111001001010110010",
						 "000101111001001110000001",
						 "000101111001010001010000",
						 "000101111001010100011111",
						 "000101111001010111101110",
						 "000101111001011010111101",
						 "000101111001011110001100",
						 "000101111001100001011011",
						 "000101111001100100101010",
						 "000101111001100111111001",
						 "000101111011011010010110",
						 "000101111011011101100101",
						 "000101111011100000110100",
						 "000101111011100100000011",
						 "000101111011100111010010",
						 "000101111011101010100001",
						 "000101111011101101110000",
						 "000101111011110000111111",
						 "000101111011110100001110",
						 "000101111011110111011101",
						 "000101111011111010101100",
						 "000101111011111101111011",
						 "000101111100000001001010",
						 "000101111100000100011001",
						 "000101111100000111101000",
						 "000101111100001010110111",
						 "000101111011011010010110",
						 "000101111011011101100101",
						 "000101111011100000110100",
						 "000101111011100100000011",
						 "000101111011100111010010",
						 "000101111011101010100001",
						 "000101111011101101110000",
						 "000101111011110000111111",
						 "000101111011110100001110",
						 "000101111011110111011101",
						 "000101111011111010101100",
						 "000101111011111101111011",
						 "000101111100000001001010",
						 "000101111100000100011001",
						 "000101111100000111101000",
						 "000101111100001010110111",
						 "000101111011011010010110",
						 "000101111011011101100101",
						 "000101111011100000110100",
						 "000101111011100100000011",
						 "000101111011100111010010",
						 "000101111011101010100001",
						 "000101111011101101110000",
						 "000101111011110000111111",
						 "000101111011110100001110",
						 "000101111011110111011101",
						 "000101111011111010101100",
						 "000101111011111101111011",
						 "000101111100000001001010",
						 "000101111100000100011001",
						 "000101111100000111101000",
						 "000101111100001010110111",
						 "000101111101111101010100",
						 "000101111110000000100010",
						 "000101111110000011110000",
						 "000101111110000110111110",
						 "000101111110001010001100",
						 "000101111110001101011010",
						 "000101111110010000101000",
						 "000101111110010011110110",
						 "000101111110010111000100",
						 "000101111110011010010010",
						 "000101111110011101100000",
						 "000101111110100000101110",
						 "000101111110100011111100",
						 "000101111110100111001010",
						 "000101111110101010011000",
						 "000101111110101101100110",
						 "000101111101111101010100",
						 "000101111110000000100010",
						 "000101111110000011110000",
						 "000101111110000110111110",
						 "000101111110001010001100",
						 "000101111110001101011010",
						 "000101111110010000101000",
						 "000101111110010011110110",
						 "000101111110010111000100",
						 "000101111110011010010010",
						 "000101111110011101100000",
						 "000101111110100000101110",
						 "000101111110100011111100",
						 "000101111110100111001010",
						 "000101111110101010011000",
						 "000101111110101101100110",
						 "000101111101111101010100",
						 "000101111110000000100010",
						 "000101111110000011110000",
						 "000101111110000110111110",
						 "000101111110001010001100",
						 "000101111110001101011010",
						 "000101111110010000101000",
						 "000101111110010011110110",
						 "000101111110010111000100",
						 "000101111110011010010010",
						 "000101111110011101100000",
						 "000101111110100000101110",
						 "000101111110100011111100",
						 "000101111110100111001010",
						 "000101111110101010011000",
						 "000101111110101101100110",
						 "000110000000100000010010",
						 "000110000000100011100000",
						 "000110000000100110101110",
						 "000110000000101001111100",
						 "000110000000101101001010",
						 "000110000000110000011000",
						 "000110000000110011100110",
						 "000110000000110110110100",
						 "000110000000111010000010",
						 "000110000000111101010000",
						 "000110000001000000011110",
						 "000110000001000011101100",
						 "000110000001000110111010",
						 "000110000001001010001000",
						 "000110000001001101010110",
						 "000110000001010000100100",
						 "000110000000100000010010",
						 "000110000000100011011111",
						 "000110000000100110101100",
						 "000110000000101001111001",
						 "000110000000101101000110",
						 "000110000000110000010011",
						 "000110000000110011100000",
						 "000110000000110110101101",
						 "000110000000111001111010",
						 "000110000000111101000111",
						 "000110000001000000010100",
						 "000110000001000011100001",
						 "000110000001000110101110",
						 "000110000001001001111011",
						 "000110000001001101001000",
						 "000110000001010000010101",
						 "000110000000100000010010",
						 "000110000000100011011111",
						 "000110000000100110101100",
						 "000110000000101001111001",
						 "000110000000101101000110",
						 "000110000000110000010011",
						 "000110000000110011100000",
						 "000110000000110110101101",
						 "000110000000111001111010",
						 "000110000000111101000111",
						 "000110000001000000010100",
						 "000110000001000011100001",
						 "000110000001000110101110",
						 "000110000001001001111011",
						 "000110000001001101001000",
						 "000110000001010000010101",
						 "000110000011000011010000",
						 "000110000011000110011101",
						 "000110000011001001101010",
						 "000110000011001100110111",
						 "000110000011010000000100",
						 "000110000011010011010001",
						 "000110000011010110011110",
						 "000110000011011001101011",
						 "000110000011011100111000",
						 "000110000011100000000101",
						 "000110000011100011010010",
						 "000110000011100110011111",
						 "000110000011101001101100",
						 "000110000011101100111001",
						 "000110000011110000000110",
						 "000110000011110011010011",
						 "000110000011000011010000",
						 "000110000011000110011101",
						 "000110000011001001101010",
						 "000110000011001100110111",
						 "000110000011010000000100",
						 "000110000011010011010001",
						 "000110000011010110011110",
						 "000110000011011001101011",
						 "000110000011011100111000",
						 "000110000011100000000101",
						 "000110000011100011010010",
						 "000110000011100110011111",
						 "000110000011101001101100",
						 "000110000011101100111001",
						 "000110000011110000000110",
						 "000110000011110011010011",
						 "000110000011000011010000",
						 "000110000011000110011100",
						 "000110000011001001101000",
						 "000110000011001100110100",
						 "000110000011010000000000",
						 "000110000011010011001100",
						 "000110000011010110011000",
						 "000110000011011001100100",
						 "000110000011011100110000",
						 "000110000011011111111100",
						 "000110000011100011001000",
						 "000110000011100110010100",
						 "000110000011101001100000",
						 "000110000011101100101100",
						 "000110000011101111111000",
						 "000110000011110011000100",
						 "000110000101100110001110",
						 "000110000101101001011010",
						 "000110000101101100100110",
						 "000110000101101111110010",
						 "000110000101110010111110",
						 "000110000101110110001010",
						 "000110000101111001010110",
						 "000110000101111100100010",
						 "000110000101111111101110",
						 "000110000110000010111010",
						 "000110000110000110000110",
						 "000110000110001001010010",
						 "000110000110001100011110",
						 "000110000110001111101010",
						 "000110000110010010110110",
						 "000110000110010110000010",
						 "000110000101100110001110",
						 "000110000101101001011010",
						 "000110000101101100100110",
						 "000110000101101111110010",
						 "000110000101110010111110",
						 "000110000101110110001010",
						 "000110000101111001010110",
						 "000110000101111100100010",
						 "000110000101111111101110",
						 "000110000110000010111010",
						 "000110000110000110000110",
						 "000110000110001001010010",
						 "000110000110001100011110",
						 "000110000110001111101010",
						 "000110000110010010110110",
						 "000110000110010110000010",
						 "000110000101100110001110",
						 "000110000101101001011010",
						 "000110000101101100100110",
						 "000110000101101111110010",
						 "000110000101110010111110",
						 "000110000101110110001010",
						 "000110000101111001010110",
						 "000110000101111100100010",
						 "000110000101111111101110",
						 "000110000110000010111010",
						 "000110000110000110000110",
						 "000110000110001001010010",
						 "000110000110001100011110",
						 "000110000110001111101010",
						 "000110000110010010110110",
						 "000110000110010110000010",
						 "000110000101100110001110",
						 "000110000101101001011010",
						 "000110000101101100100110",
						 "000110000101101111110010",
						 "000110000101110010111110",
						 "000110000101110110001010",
						 "000110000101111001010110",
						 "000110000101111100100010",
						 "000110000101111111101110",
						 "000110000110000010111010",
						 "000110000110000110000110",
						 "000110000110001001010010",
						 "000110000110001100011110",
						 "000110000110001111101010",
						 "000110000110010010110110",
						 "000110000110010110000010",
						 "000110001000001001001100",
						 "000110001000001100010111",
						 "000110001000001111100010",
						 "000110001000010010101101",
						 "000110001000010101111000",
						 "000110001000011001000011",
						 "000110001000011100001110",
						 "000110001000011111011001",
						 "000110001000100010100100",
						 "000110001000100101101111",
						 "000110001000101000111010",
						 "000110001000101100000101",
						 "000110001000101111010000",
						 "000110001000110010011011",
						 "000110001000110101100110",
						 "000110001000111000110001",
						 "000110001000001001001100",
						 "000110001000001100010111",
						 "000110001000001111100010",
						 "000110001000010010101101",
						 "000110001000010101111000",
						 "000110001000011001000011",
						 "000110001000011100001110",
						 "000110001000011111011001",
						 "000110001000100010100100",
						 "000110001000100101101111",
						 "000110001000101000111010",
						 "000110001000101100000101",
						 "000110001000101111010000",
						 "000110001000110010011011",
						 "000110001000110101100110",
						 "000110001000111000110001",
						 "000110001000001001001100",
						 "000110001000001100010111",
						 "000110001000001111100010",
						 "000110001000010010101101",
						 "000110001000010101111000",
						 "000110001000011001000011",
						 "000110001000011100001110",
						 "000110001000011111011001",
						 "000110001000100010100100",
						 "000110001000100101101111",
						 "000110001000101000111010",
						 "000110001000101100000101",
						 "000110001000101111010000",
						 "000110001000110010011011",
						 "000110001000110101100110",
						 "000110001000111000110001",
						 "000110001010101100001010",
						 "000110001010101111010101",
						 "000110001010110010100000",
						 "000110001010110101101011",
						 "000110001010111000110110",
						 "000110001010111100000001",
						 "000110001010111111001100",
						 "000110001011000010010111",
						 "000110001011000101100010",
						 "000110001011001000101101",
						 "000110001011001011111000",
						 "000110001011001111000011",
						 "000110001011010010001110",
						 "000110001011010101011001",
						 "000110001011011000100100",
						 "000110001011011011101111",
						 "000110001010101100001010",
						 "000110001010101111010100",
						 "000110001010110010011110",
						 "000110001010110101101000",
						 "000110001010111000110010",
						 "000110001010111011111100",
						 "000110001010111111000110",
						 "000110001011000010010000",
						 "000110001011000101011010",
						 "000110001011001000100100",
						 "000110001011001011101110",
						 "000110001011001110111000",
						 "000110001011010010000010",
						 "000110001011010101001100",
						 "000110001011011000010110",
						 "000110001011011011100000",
						 "000110001010101100001010",
						 "000110001010101111010100",
						 "000110001010110010011110",
						 "000110001010110101101000",
						 "000110001010111000110010",
						 "000110001010111011111100",
						 "000110001010111111000110",
						 "000110001011000010010000",
						 "000110001011000101011010",
						 "000110001011001000100100",
						 "000110001011001011101110",
						 "000110001011001110111000",
						 "000110001011010010000010",
						 "000110001011010101001100",
						 "000110001011011000010110",
						 "000110001011011011100000",
						 "000110001101001111001000",
						 "000110001101010010010010",
						 "000110001101010101011100",
						 "000110001101011000100110",
						 "000110001101011011110000",
						 "000110001101011110111010",
						 "000110001101100010000100",
						 "000110001101100101001110",
						 "000110001101101000011000",
						 "000110001101101011100010",
						 "000110001101101110101100",
						 "000110001101110001110110",
						 "000110001101110101000000",
						 "000110001101111000001010",
						 "000110001101111011010100",
						 "000110001101111110011110",
						 "000110001101001111001000",
						 "000110001101010010010010",
						 "000110001101010101011100",
						 "000110001101011000100110",
						 "000110001101011011110000",
						 "000110001101011110111010",
						 "000110001101100010000100",
						 "000110001101100101001110",
						 "000110001101101000011000",
						 "000110001101101011100010",
						 "000110001101101110101100",
						 "000110001101110001110110",
						 "000110001101110101000000",
						 "000110001101111000001010",
						 "000110001101111011010100",
						 "000110001101111110011110",
						 "000110001101001111001000",
						 "000110001101010010010001",
						 "000110001101010101011010",
						 "000110001101011000100011",
						 "000110001101011011101100",
						 "000110001101011110110101",
						 "000110001101100001111110",
						 "000110001101100101000111",
						 "000110001101101000010000",
						 "000110001101101011011001",
						 "000110001101101110100010",
						 "000110001101110001101011",
						 "000110001101110100110100",
						 "000110001101110111111101",
						 "000110001101111011000110",
						 "000110001101111110001111",
						 "000110001111110010000110",
						 "000110001111110101001111",
						 "000110001111111000011000",
						 "000110001111111011100001",
						 "000110001111111110101010",
						 "000110010000000001110011",
						 "000110010000000100111100",
						 "000110010000001000000101",
						 "000110010000001011001110",
						 "000110010000001110010111",
						 "000110010000010001100000",
						 "000110010000010100101001",
						 "000110010000010111110010",
						 "000110010000011010111011",
						 "000110010000011110000100",
						 "000110010000100001001101",
						 "000110001111110010000110",
						 "000110001111110101001111",
						 "000110001111111000011000",
						 "000110001111111011100001",
						 "000110001111111110101010",
						 "000110010000000001110011",
						 "000110010000000100111100",
						 "000110010000001000000101",
						 "000110010000001011001110",
						 "000110010000001110010111",
						 "000110010000010001100000",
						 "000110010000010100101001",
						 "000110010000010111110010",
						 "000110010000011010111011",
						 "000110010000011110000100",
						 "000110010000100001001101",
						 "000110001111110010000110",
						 "000110001111110101001111",
						 "000110001111111000011000",
						 "000110001111111011100001",
						 "000110001111111110101010",
						 "000110010000000001110011",
						 "000110010000000100111100",
						 "000110010000001000000101",
						 "000110010000001011001110",
						 "000110010000001110010111",
						 "000110010000010001100000",
						 "000110010000010100101001",
						 "000110010000010111110010",
						 "000110010000011010111011",
						 "000110010000011110000100",
						 "000110010000100001001101",
						 "000110010010010101000100",
						 "000110010010011000001100",
						 "000110010010011011010100",
						 "000110010010011110011100",
						 "000110010010100001100100",
						 "000110010010100100101100",
						 "000110010010100111110100",
						 "000110010010101010111100",
						 "000110010010101110000100",
						 "000110010010110001001100",
						 "000110010010110100010100",
						 "000110010010110111011100",
						 "000110010010111010100100",
						 "000110010010111101101100",
						 "000110010011000000110100",
						 "000110010011000011111100",
						 "000110010010010101000100",
						 "000110010010011000001100",
						 "000110010010011011010100",
						 "000110010010011110011100",
						 "000110010010100001100100",
						 "000110010010100100101100",
						 "000110010010100111110100",
						 "000110010010101010111100",
						 "000110010010101110000100",
						 "000110010010110001001100",
						 "000110010010110100010100",
						 "000110010010110111011100",
						 "000110010010111010100100",
						 "000110010010111101101100",
						 "000110010011000000110100",
						 "000110010011000011111100",
						 "000110010010010101000100",
						 "000110010010011000001100",
						 "000110010010011011010100",
						 "000110010010011110011100",
						 "000110010010100001100100",
						 "000110010010100100101100",
						 "000110010010100111110100",
						 "000110010010101010111100",
						 "000110010010101110000100",
						 "000110010010110001001100",
						 "000110010010110100010100",
						 "000110010010110111011100",
						 "000110010010111010100100",
						 "000110010010111101101100",
						 "000110010011000000110100",
						 "000110010011000011111100",
						 "000110010010010101000100",
						 "000110010010011000001100",
						 "000110010010011011010100",
						 "000110010010011110011100",
						 "000110010010100001100100",
						 "000110010010100100101100",
						 "000110010010100111110100",
						 "000110010010101010111100",
						 "000110010010101110000100",
						 "000110010010110001001100",
						 "000110010010110100010100",
						 "000110010010110111011100",
						 "000110010010111010100100",
						 "000110010010111101101100",
						 "000110010011000000110100",
						 "000110010011000011111100",
						 "000110010100111000000010",
						 "000110010100111011001001",
						 "000110010100111110010000",
						 "000110010101000001010111",
						 "000110010101000100011110",
						 "000110010101000111100101",
						 "000110010101001010101100",
						 "000110010101001101110011",
						 "000110010101010000111010",
						 "000110010101010100000001",
						 "000110010101010111001000",
						 "000110010101011010001111",
						 "000110010101011101010110",
						 "000110010101100000011101",
						 "000110010101100011100100",
						 "000110010101100110101011",
						 "000110010100111000000010",
						 "000110010100111011001001",
						 "000110010100111110010000",
						 "000110010101000001010111",
						 "000110010101000100011110",
						 "000110010101000111100101",
						 "000110010101001010101100",
						 "000110010101001101110011",
						 "000110010101010000111010",
						 "000110010101010100000001",
						 "000110010101010111001000",
						 "000110010101011010001111",
						 "000110010101011101010110",
						 "000110010101100000011101",
						 "000110010101100011100100",
						 "000110010101100110101011",
						 "000110010100111000000010",
						 "000110010100111011001001",
						 "000110010100111110010000",
						 "000110010101000001010111",
						 "000110010101000100011110",
						 "000110010101000111100101",
						 "000110010101001010101100",
						 "000110010101001101110011",
						 "000110010101010000111010",
						 "000110010101010100000001",
						 "000110010101010111001000",
						 "000110010101011010001111",
						 "000110010101011101010110",
						 "000110010101100000011101",
						 "000110010101100011100100",
						 "000110010101100110101011",
						 "000110010111011011000000",
						 "000110010111011110000111",
						 "000110010111100001001110",
						 "000110010111100100010101",
						 "000110010111100111011100",
						 "000110010111101010100011",
						 "000110010111101101101010",
						 "000110010111110000110001",
						 "000110010111110011111000",
						 "000110010111110110111111",
						 "000110010111111010000110",
						 "000110010111111101001101",
						 "000110011000000000010100",
						 "000110011000000011011011",
						 "000110011000000110100010",
						 "000110011000001001101001",
						 "000110010111011011000000",
						 "000110010111011110000110",
						 "000110010111100001001100",
						 "000110010111100100010010",
						 "000110010111100111011000",
						 "000110010111101010011110",
						 "000110010111101101100100",
						 "000110010111110000101010",
						 "000110010111110011110000",
						 "000110010111110110110110",
						 "000110010111111001111100",
						 "000110010111111101000010",
						 "000110011000000000001000",
						 "000110011000000011001110",
						 "000110011000000110010100",
						 "000110011000001001011010",
						 "000110010111011011000000",
						 "000110010111011110000110",
						 "000110010111100001001100",
						 "000110010111100100010010",
						 "000110010111100111011000",
						 "000110010111101010011110",
						 "000110010111101101100100",
						 "000110010111110000101010",
						 "000110010111110011110000",
						 "000110010111110110110110",
						 "000110010111111001111100",
						 "000110010111111101000010",
						 "000110011000000000001000",
						 "000110011000000011001110",
						 "000110011000000110010100",
						 "000110011000001001011010",
						 "000110011001111101111110",
						 "000110011010000001000100",
						 "000110011010000100001010",
						 "000110011010000111010000",
						 "000110011010001010010110",
						 "000110011010001101011100",
						 "000110011010010000100010",
						 "000110011010010011101000",
						 "000110011010010110101110",
						 "000110011010011001110100",
						 "000110011010011100111010",
						 "000110011010100000000000",
						 "000110011010100011000110",
						 "000110011010100110001100",
						 "000110011010101001010010",
						 "000110011010101100011000",
						 "000110011001111101111110",
						 "000110011010000001000100",
						 "000110011010000100001010",
						 "000110011010000111010000",
						 "000110011010001010010110",
						 "000110011010001101011100",
						 "000110011010010000100010",
						 "000110011010010011101000",
						 "000110011010010110101110",
						 "000110011010011001110100",
						 "000110011010011100111010",
						 "000110011010100000000000",
						 "000110011010100011000110",
						 "000110011010100110001100",
						 "000110011010101001010010",
						 "000110011010101100011000",
						 "000110011001111101111110",
						 "000110011010000001000011",
						 "000110011010000100001000",
						 "000110011010000111001101",
						 "000110011010001010010010",
						 "000110011010001101010111",
						 "000110011010010000011100",
						 "000110011010010011100001",
						 "000110011010010110100110",
						 "000110011010011001101011",
						 "000110011010011100110000",
						 "000110011010011111110101",
						 "000110011010100010111010",
						 "000110011010100101111111",
						 "000110011010101001000100",
						 "000110011010101100001001",
						 "000110011001111101111110",
						 "000110011010000001000011",
						 "000110011010000100001000",
						 "000110011010000111001101",
						 "000110011010001010010010",
						 "000110011010001101010111",
						 "000110011010010000011100",
						 "000110011010010011100001",
						 "000110011010010110100110",
						 "000110011010011001101011",
						 "000110011010011100110000",
						 "000110011010011111110101",
						 "000110011010100010111010",
						 "000110011010100101111111",
						 "000110011010101001000100",
						 "000110011010101100001001",
						 "000110011100100000111100",
						 "000110011100100100000001",
						 "000110011100100111000110",
						 "000110011100101010001011",
						 "000110011100101101010000",
						 "000110011100110000010101",
						 "000110011100110011011010",
						 "000110011100110110011111",
						 "000110011100111001100100",
						 "000110011100111100101001",
						 "000110011100111111101110",
						 "000110011101000010110011",
						 "000110011101000101111000",
						 "000110011101001000111101",
						 "000110011101001100000010",
						 "000110011101001111000111",
						 "000110011100100000111100",
						 "000110011100100100000001",
						 "000110011100100111000110",
						 "000110011100101010001011",
						 "000110011100101101010000",
						 "000110011100110000010101",
						 "000110011100110011011010",
						 "000110011100110110011111",
						 "000110011100111001100100",
						 "000110011100111100101001",
						 "000110011100111111101110",
						 "000110011101000010110011",
						 "000110011101000101111000",
						 "000110011101001000111101",
						 "000110011101001100000010",
						 "000110011101001111000111",
						 "000110011100100000111100",
						 "000110011100100100000000",
						 "000110011100100111000100",
						 "000110011100101010001000",
						 "000110011100101101001100",
						 "000110011100110000010000",
						 "000110011100110011010100",
						 "000110011100110110011000",
						 "000110011100111001011100",
						 "000110011100111100100000",
						 "000110011100111111100100",
						 "000110011101000010101000",
						 "000110011101000101101100",
						 "000110011101001000110000",
						 "000110011101001011110100",
						 "000110011101001110111000",
						 "000110011111000011111010",
						 "000110011111000110111110",
						 "000110011111001010000010",
						 "000110011111001101000110",
						 "000110011111010000001010",
						 "000110011111010011001110",
						 "000110011111010110010010",
						 "000110011111011001010110",
						 "000110011111011100011010",
						 "000110011111011111011110",
						 "000110011111100010100010",
						 "000110011111100101100110",
						 "000110011111101000101010",
						 "000110011111101011101110",
						 "000110011111101110110010",
						 "000110011111110001110110",
						 "000110011111000011111010",
						 "000110011111000110111110",
						 "000110011111001010000010",
						 "000110011111001101000110",
						 "000110011111010000001010",
						 "000110011111010011001110",
						 "000110011111010110010010",
						 "000110011111011001010110",
						 "000110011111011100011010",
						 "000110011111011111011110",
						 "000110011111100010100010",
						 "000110011111100101100110",
						 "000110011111101000101010",
						 "000110011111101011101110",
						 "000110011111101110110010",
						 "000110011111110001110110",
						 "000110011111000011111010",
						 "000110011111000110111110",
						 "000110011111001010000010",
						 "000110011111001101000110",
						 "000110011111010000001010",
						 "000110011111010011001110",
						 "000110011111010110010010",
						 "000110011111011001010110",
						 "000110011111011100011010",
						 "000110011111011111011110",
						 "000110011111100010100010",
						 "000110011111100101100110",
						 "000110011111101000101010",
						 "000110011111101011101110",
						 "000110011111101110110010",
						 "000110011111110001110110",
						 "000110100001100110111000",
						 "000110100001101001111011",
						 "000110100001101100111110",
						 "000110100001110000000001",
						 "000110100001110011000100",
						 "000110100001110110000111",
						 "000110100001111001001010",
						 "000110100001111100001101",
						 "000110100001111111010000",
						 "000110100010000010010011",
						 "000110100010000101010110",
						 "000110100010001000011001",
						 "000110100010001011011100",
						 "000110100010001110011111",
						 "000110100010010001100010",
						 "000110100010010100100101",
						 "000110100001100110111000",
						 "000110100001101001111011",
						 "000110100001101100111110",
						 "000110100001110000000001",
						 "000110100001110011000100",
						 "000110100001110110000111",
						 "000110100001111001001010",
						 "000110100001111100001101",
						 "000110100001111111010000",
						 "000110100010000010010011",
						 "000110100010000101010110",
						 "000110100010001000011001",
						 "000110100010001011011100",
						 "000110100010001110011111",
						 "000110100010010001100010",
						 "000110100010010100100101",
						 "000110100001100110111000",
						 "000110100001101001111011",
						 "000110100001101100111110",
						 "000110100001110000000001",
						 "000110100001110011000100",
						 "000110100001110110000111",
						 "000110100001111001001010",
						 "000110100001111100001101",
						 "000110100001111111010000",
						 "000110100010000010010011",
						 "000110100010000101010110",
						 "000110100010001000011001",
						 "000110100010001011011100",
						 "000110100010001110011111",
						 "000110100010010001100010",
						 "000110100010010100100101",
						 "000110100001100110111000",
						 "000110100001101001111011",
						 "000110100001101100111110",
						 "000110100001110000000001",
						 "000110100001110011000100",
						 "000110100001110110000111",
						 "000110100001111001001010",
						 "000110100001111100001101",
						 "000110100001111111010000",
						 "000110100010000010010011",
						 "000110100010000101010110",
						 "000110100010001000011001",
						 "000110100010001011011100",
						 "000110100010001110011111",
						 "000110100010010001100010",
						 "000110100010010100100101",
						 "000110100100001001110110",
						 "000110100100001100111000",
						 "000110100100001111111010",
						 "000110100100010010111100",
						 "000110100100010101111110",
						 "000110100100011001000000",
						 "000110100100011100000010",
						 "000110100100011111000100",
						 "000110100100100010000110",
						 "000110100100100101001000",
						 "000110100100101000001010",
						 "000110100100101011001100",
						 "000110100100101110001110",
						 "000110100100110001010000",
						 "000110100100110100010010",
						 "000110100100110111010100",
						 "000110100100001001110110",
						 "000110100100001100111000",
						 "000110100100001111111010",
						 "000110100100010010111100",
						 "000110100100010101111110",
						 "000110100100011001000000",
						 "000110100100011100000010",
						 "000110100100011111000100",
						 "000110100100100010000110",
						 "000110100100100101001000",
						 "000110100100101000001010",
						 "000110100100101011001100",
						 "000110100100101110001110",
						 "000110100100110001010000",
						 "000110100100110100010010",
						 "000110100100110111010100",
						 "000110100100001001110110",
						 "000110100100001100111000",
						 "000110100100001111111010",
						 "000110100100010010111100",
						 "000110100100010101111110",
						 "000110100100011001000000",
						 "000110100100011100000010",
						 "000110100100011111000100",
						 "000110100100100010000110",
						 "000110100100100101001000",
						 "000110100100101000001010",
						 "000110100100101011001100",
						 "000110100100101110001110",
						 "000110100100110001010000",
						 "000110100100110100010010",
						 "000110100100110111010100",
						 "000110100110101100110100",
						 "000110100110101111110110",
						 "000110100110110010111000",
						 "000110100110110101111010",
						 "000110100110111000111100",
						 "000110100110111011111110",
						 "000110100110111111000000",
						 "000110100111000010000010",
						 "000110100111000101000100",
						 "000110100111001000000110",
						 "000110100111001011001000",
						 "000110100111001110001010",
						 "000110100111010001001100",
						 "000110100111010100001110",
						 "000110100111010111010000",
						 "000110100111011010010010",
						 "000110100110101100110100",
						 "000110100110101111110101",
						 "000110100110110010110110",
						 "000110100110110101110111",
						 "000110100110111000111000",
						 "000110100110111011111001",
						 "000110100110111110111010",
						 "000110100111000001111011",
						 "000110100111000100111100",
						 "000110100111000111111101",
						 "000110100111001010111110",
						 "000110100111001101111111",
						 "000110100111010001000000",
						 "000110100111010100000001",
						 "000110100111010111000010",
						 "000110100111011010000011",
						 "000110100110101100110100",
						 "000110100110101111110101",
						 "000110100110110010110110",
						 "000110100110110101110111",
						 "000110100110111000111000",
						 "000110100110111011111001",
						 "000110100110111110111010",
						 "000110100111000001111011",
						 "000110100111000100111100",
						 "000110100111000111111101",
						 "000110100111001010111110",
						 "000110100111001101111111",
						 "000110100111010001000000",
						 "000110100111010100000001",
						 "000110100111010111000010",
						 "000110100111011010000011",
						 "000110101001001111110010",
						 "000110101001010010110011",
						 "000110101001010101110100",
						 "000110101001011000110101",
						 "000110101001011011110110",
						 "000110101001011110110111",
						 "000110101001100001111000",
						 "000110101001100100111001",
						 "000110101001100111111010",
						 "000110101001101010111011",
						 "000110101001101101111100",
						 "000110101001110000111101",
						 "000110101001110011111110",
						 "000110101001110110111111",
						 "000110101001111010000000",
						 "000110101001111101000001",
						 "000110101001001111110010",
						 "000110101001010010110011",
						 "000110101001010101110100",
						 "000110101001011000110101",
						 "000110101001011011110110",
						 "000110101001011110110111",
						 "000110101001100001111000",
						 "000110101001100100111001",
						 "000110101001100111111010",
						 "000110101001101010111011",
						 "000110101001101101111100",
						 "000110101001110000111101",
						 "000110101001110011111110",
						 "000110101001110110111111",
						 "000110101001111010000000",
						 "000110101001111101000001",
						 "000110101001001111110010",
						 "000110101001010010110010",
						 "000110101001010101110010",
						 "000110101001011000110010",
						 "000110101001011011110010",
						 "000110101001011110110010",
						 "000110101001100001110010",
						 "000110101001100100110010",
						 "000110101001100111110010",
						 "000110101001101010110010",
						 "000110101001101101110010",
						 "000110101001110000110010",
						 "000110101001110011110010",
						 "000110101001110110110010",
						 "000110101001111001110010",
						 "000110101001111100110010",
						 "000110101001001111110010",
						 "000110101001010010110010",
						 "000110101001010101110010",
						 "000110101001011000110010",
						 "000110101001011011110010",
						 "000110101001011110110010",
						 "000110101001100001110010",
						 "000110101001100100110010",
						 "000110101001100111110010",
						 "000110101001101010110010",
						 "000110101001101101110010",
						 "000110101001110000110010",
						 "000110101001110011110010",
						 "000110101001110110110010",
						 "000110101001111001110010",
						 "000110101001111100110010",
						 "000110101011110010110000",
						 "000110101011110101110000",
						 "000110101011111000110000",
						 "000110101011111011110000",
						 "000110101011111110110000",
						 "000110101100000001110000",
						 "000110101100000100110000",
						 "000110101100000111110000",
						 "000110101100001010110000",
						 "000110101100001101110000",
						 "000110101100010000110000",
						 "000110101100010011110000",
						 "000110101100010110110000",
						 "000110101100011001110000",
						 "000110101100011100110000",
						 "000110101100011111110000",
						 "000110101011110010110000",
						 "000110101011110101110000",
						 "000110101011111000110000",
						 "000110101011111011110000",
						 "000110101011111110110000",
						 "000110101100000001110000",
						 "000110101100000100110000",
						 "000110101100000111110000",
						 "000110101100001010110000",
						 "000110101100001101110000",
						 "000110101100010000110000",
						 "000110101100010011110000",
						 "000110101100010110110000",
						 "000110101100011001110000",
						 "000110101100011100110000",
						 "000110101100011111110000",
						 "000110101011110010110000",
						 "000110101011110101101111",
						 "000110101011111000101110",
						 "000110101011111011101101",
						 "000110101011111110101100",
						 "000110101100000001101011",
						 "000110101100000100101010",
						 "000110101100000111101001",
						 "000110101100001010101000",
						 "000110101100001101100111",
						 "000110101100010000100110",
						 "000110101100010011100101",
						 "000110101100010110100100",
						 "000110101100011001100011",
						 "000110101100011100100010",
						 "000110101100011111100001",
						 "000110101110010101101110",
						 "000110101110011000101101",
						 "000110101110011011101100",
						 "000110101110011110101011",
						 "000110101110100001101010",
						 "000110101110100100101001",
						 "000110101110100111101000",
						 "000110101110101010100111",
						 "000110101110101101100110",
						 "000110101110110000100101",
						 "000110101110110011100100",
						 "000110101110110110100011",
						 "000110101110111001100010",
						 "000110101110111100100001",
						 "000110101110111111100000",
						 "000110101111000010011111",
						 "000110101110010101101110",
						 "000110101110011000101101",
						 "000110101110011011101100",
						 "000110101110011110101011",
						 "000110101110100001101010",
						 "000110101110100100101001",
						 "000110101110100111101000",
						 "000110101110101010100111",
						 "000110101110101101100110",
						 "000110101110110000100101",
						 "000110101110110011100100",
						 "000110101110110110100011",
						 "000110101110111001100010",
						 "000110101110111100100001",
						 "000110101110111111100000",
						 "000110101111000010011111",
						 "000110101110010101101110",
						 "000110101110011000101101",
						 "000110101110011011101100",
						 "000110101110011110101011",
						 "000110101110100001101010",
						 "000110101110100100101001",
						 "000110101110100111101000",
						 "000110101110101010100111",
						 "000110101110101101100110",
						 "000110101110110000100101",
						 "000110101110110011100100",
						 "000110101110110110100011",
						 "000110101110111001100010",
						 "000110101110111100100001",
						 "000110101110111111100000",
						 "000110101111000010011111",
						 "000110110000111000101100",
						 "000110110000111011101010",
						 "000110110000111110101000",
						 "000110110001000001100110",
						 "000110110001000100100100",
						 "000110110001000111100010",
						 "000110110001001010100000",
						 "000110110001001101011110",
						 "000110110001010000011100",
						 "000110110001010011011010",
						 "000110110001010110011000",
						 "000110110001011001010110",
						 "000110110001011100010100",
						 "000110110001011111010010",
						 "000110110001100010010000",
						 "000110110001100101001110",
						 "000110110000111000101100",
						 "000110110000111011101010",
						 "000110110000111110101000",
						 "000110110001000001100110",
						 "000110110001000100100100",
						 "000110110001000111100010",
						 "000110110001001010100000",
						 "000110110001001101011110",
						 "000110110001010000011100",
						 "000110110001010011011010",
						 "000110110001010110011000",
						 "000110110001011001010110",
						 "000110110001011100010100",
						 "000110110001011111010010",
						 "000110110001100010010000",
						 "000110110001100101001110",
						 "000110110000111000101100",
						 "000110110000111011101010",
						 "000110110000111110101000",
						 "000110110001000001100110",
						 "000110110001000100100100",
						 "000110110001000111100010",
						 "000110110001001010100000",
						 "000110110001001101011110",
						 "000110110001010000011100",
						 "000110110001010011011010",
						 "000110110001010110011000",
						 "000110110001011001010110",
						 "000110110001011100010100",
						 "000110110001011111010010",
						 "000110110001100010010000",
						 "000110110001100101001110",
						 "000110110000111000101100",
						 "000110110000111011101010",
						 "000110110000111110101000",
						 "000110110001000001100110",
						 "000110110001000100100100",
						 "000110110001000111100010",
						 "000110110001001010100000",
						 "000110110001001101011110",
						 "000110110001010000011100",
						 "000110110001010011011010",
						 "000110110001010110011000",
						 "000110110001011001010110",
						 "000110110001011100010100",
						 "000110110001011111010010",
						 "000110110001100010010000",
						 "000110110001100101001110",
						 "000110110011011011101010",
						 "000110110011011110100111",
						 "000110110011100001100100",
						 "000110110011100100100001",
						 "000110110011100111011110",
						 "000110110011101010011011",
						 "000110110011101101011000",
						 "000110110011110000010101",
						 "000110110011110011010010",
						 "000110110011110110001111",
						 "000110110011111001001100",
						 "000110110011111100001001",
						 "000110110011111111000110",
						 "000110110100000010000011",
						 "000110110100000101000000",
						 "000110110100000111111101",
						 "000110110011011011101010",
						 "000110110011011110100111",
						 "000110110011100001100100",
						 "000110110011100100100001",
						 "000110110011100111011110",
						 "000110110011101010011011",
						 "000110110011101101011000",
						 "000110110011110000010101",
						 "000110110011110011010010",
						 "000110110011110110001111",
						 "000110110011111001001100",
						 "000110110011111100001001",
						 "000110110011111111000110",
						 "000110110100000010000011",
						 "000110110100000101000000",
						 "000110110100000111111101",
						 "000110110011011011101010",
						 "000110110011011110100111",
						 "000110110011100001100100",
						 "000110110011100100100001",
						 "000110110011100111011110",
						 "000110110011101010011011",
						 "000110110011101101011000",
						 "000110110011110000010101",
						 "000110110011110011010010",
						 "000110110011110110001111",
						 "000110110011111001001100",
						 "000110110011111100001001",
						 "000110110011111111000110",
						 "000110110100000010000011",
						 "000110110100000101000000",
						 "000110110100000111111101",
						 "000110110101111110101000",
						 "000110110110000001100101",
						 "000110110110000100100010",
						 "000110110110000111011111",
						 "000110110110001010011100",
						 "000110110110001101011001",
						 "000110110110010000010110",
						 "000110110110010011010011",
						 "000110110110010110010000",
						 "000110110110011001001101",
						 "000110110110011100001010",
						 "000110110110011111000111",
						 "000110110110100010000100",
						 "000110110110100101000001",
						 "000110110110100111111110",
						 "000110110110101010111011",
						 "000110110101111110101000",
						 "000110110110000001100100",
						 "000110110110000100100000",
						 "000110110110000111011100",
						 "000110110110001010011000",
						 "000110110110001101010100",
						 "000110110110010000010000",
						 "000110110110010011001100",
						 "000110110110010110001000",
						 "000110110110011001000100",
						 "000110110110011100000000",
						 "000110110110011110111100",
						 "000110110110100001111000",
						 "000110110110100100110100",
						 "000110110110100111110000",
						 "000110110110101010101100",
						 "000110110101111110101000",
						 "000110110110000001100100",
						 "000110110110000100100000",
						 "000110110110000111011100",
						 "000110110110001010011000",
						 "000110110110001101010100",
						 "000110110110010000010000",
						 "000110110110010011001100",
						 "000110110110010110001000",
						 "000110110110011001000100",
						 "000110110110011100000000",
						 "000110110110011110111100",
						 "000110110110100001111000",
						 "000110110110100100110100",
						 "000110110110100111110000",
						 "000110110110101010101100",
						 "000110110101111110101000",
						 "000110110110000001100100",
						 "000110110110000100100000",
						 "000110110110000111011100",
						 "000110110110001010011000",
						 "000110110110001101010100",
						 "000110110110010000010000",
						 "000110110110010011001100",
						 "000110110110010110001000",
						 "000110110110011001000100",
						 "000110110110011100000000",
						 "000110110110011110111100",
						 "000110110110100001111000",
						 "000110110110100100110100",
						 "000110110110100111110000",
						 "000110110110101010101100",
						 "000110111000100001100110",
						 "000110111000100100100001",
						 "000110111000100111011100",
						 "000110111000101010010111",
						 "000110111000101101010010",
						 "000110111000110000001101",
						 "000110111000110011001000",
						 "000110111000110110000011",
						 "000110111000111000111110",
						 "000110111000111011111001",
						 "000110111000111110110100",
						 "000110111001000001101111",
						 "000110111001000100101010",
						 "000110111001000111100101",
						 "000110111001001010100000",
						 "000110111001001101011011",
						 "000110111000100001100110",
						 "000110111000100100100001",
						 "000110111000100111011100",
						 "000110111000101010010111",
						 "000110111000101101010010",
						 "000110111000110000001101",
						 "000110111000110011001000",
						 "000110111000110110000011",
						 "000110111000111000111110",
						 "000110111000111011111001",
						 "000110111000111110110100",
						 "000110111001000001101111",
						 "000110111001000100101010",
						 "000110111001000111100101",
						 "000110111001001010100000",
						 "000110111001001101011011",
						 "000110111000100001100110",
						 "000110111000100100100001",
						 "000110111000100111011100",
						 "000110111000101010010111",
						 "000110111000101101010010",
						 "000110111000110000001101",
						 "000110111000110011001000",
						 "000110111000110110000011",
						 "000110111000111000111110",
						 "000110111000111011111001",
						 "000110111000111110110100",
						 "000110111001000001101111",
						 "000110111001000100101010",
						 "000110111001000111100101",
						 "000110111001001010100000",
						 "000110111001001101011011",
						 "000110111011000100100100",
						 "000110111011000111011111",
						 "000110111011001010011010",
						 "000110111011001101010101",
						 "000110111011010000010000",
						 "000110111011010011001011",
						 "000110111011010110000110",
						 "000110111011011001000001",
						 "000110111011011011111100",
						 "000110111011011110110111",
						 "000110111011100001110010",
						 "000110111011100100101101",
						 "000110111011100111101000",
						 "000110111011101010100011",
						 "000110111011101101011110",
						 "000110111011110000011001",
						 "000110111011000100100100",
						 "000110111011000111011110",
						 "000110111011001010011000",
						 "000110111011001101010010",
						 "000110111011010000001100",
						 "000110111011010011000110",
						 "000110111011010110000000",
						 "000110111011011000111010",
						 "000110111011011011110100",
						 "000110111011011110101110",
						 "000110111011100001101000",
						 "000110111011100100100010",
						 "000110111011100111011100",
						 "000110111011101010010110",
						 "000110111011101101010000",
						 "000110111011110000001010",
						 "000110111011000100100100",
						 "000110111011000111011110",
						 "000110111011001010011000",
						 "000110111011001101010010",
						 "000110111011010000001100",
						 "000110111011010011000110",
						 "000110111011010110000000",
						 "000110111011011000111010",
						 "000110111011011011110100",
						 "000110111011011110101110",
						 "000110111011100001101000",
						 "000110111011100100100010",
						 "000110111011100111011100",
						 "000110111011101010010110",
						 "000110111011101101010000",
						 "000110111011110000001010",
						 "000110111011000100100100",
						 "000110111011000111011110",
						 "000110111011001010011000",
						 "000110111011001101010010",
						 "000110111011010000001100",
						 "000110111011010011000110",
						 "000110111011010110000000",
						 "000110111011011000111010",
						 "000110111011011011110100",
						 "000110111011011110101110",
						 "000110111011100001101000",
						 "000110111011100100100010",
						 "000110111011100111011100",
						 "000110111011101010010110",
						 "000110111011101101010000",
						 "000110111011110000001010",
						 "000110111101100111100010",
						 "000110111101101010011100",
						 "000110111101101101010110",
						 "000110111101110000010000",
						 "000110111101110011001010",
						 "000110111101110110000100",
						 "000110111101111000111110",
						 "000110111101111011111000",
						 "000110111101111110110010",
						 "000110111110000001101100",
						 "000110111110000100100110",
						 "000110111110000111100000",
						 "000110111110001010011010",
						 "000110111110001101010100",
						 "000110111110010000001110",
						 "000110111110010011001000",
						 "000110111101100111100010",
						 "000110111101101010011011",
						 "000110111101101101010100",
						 "000110111101110000001101",
						 "000110111101110011000110",
						 "000110111101110101111111",
						 "000110111101111000111000",
						 "000110111101111011110001",
						 "000110111101111110101010",
						 "000110111110000001100011",
						 "000110111110000100011100",
						 "000110111110000111010101",
						 "000110111110001010001110",
						 "000110111110001101000111",
						 "000110111110010000000000",
						 "000110111110010010111001",
						 "000110111101100111100010",
						 "000110111101101010011011",
						 "000110111101101101010100",
						 "000110111101110000001101",
						 "000110111101110011000110",
						 "000110111101110101111111",
						 "000110111101111000111000",
						 "000110111101111011110001",
						 "000110111101111110101010",
						 "000110111110000001100011",
						 "000110111110000100011100",
						 "000110111110000111010101",
						 "000110111110001010001110",
						 "000110111110001101000111",
						 "000110111110010000000000",
						 "000110111110010010111001",
						 "000111000000001010100000",
						 "000111000000001101011001",
						 "000111000000010000010010",
						 "000111000000010011001011",
						 "000111000000010110000100",
						 "000111000000011000111101",
						 "000111000000011011110110",
						 "000111000000011110101111",
						 "000111000000100001101000",
						 "000111000000100100100001",
						 "000111000000100111011010",
						 "000111000000101010010011",
						 "000111000000101101001100",
						 "000111000000110000000101",
						 "000111000000110010111110",
						 "000111000000110101110111",
						 "000111000000001010100000",
						 "000111000000001101011001",
						 "000111000000010000010010",
						 "000111000000010011001011",
						 "000111000000010110000100",
						 "000111000000011000111101",
						 "000111000000011011110110",
						 "000111000000011110101111",
						 "000111000000100001101000",
						 "000111000000100100100001",
						 "000111000000100111011010",
						 "000111000000101010010011",
						 "000111000000101101001100",
						 "000111000000110000000101",
						 "000111000000110010111110",
						 "000111000000110101110111",
						 "000111000000001010100000",
						 "000111000000001101011000",
						 "000111000000010000010000",
						 "000111000000010011001000",
						 "000111000000010110000000",
						 "000111000000011000111000",
						 "000111000000011011110000",
						 "000111000000011110101000",
						 "000111000000100001100000",
						 "000111000000100100011000",
						 "000111000000100111010000",
						 "000111000000101010001000",
						 "000111000000101101000000",
						 "000111000000101111111000",
						 "000111000000110010110000",
						 "000111000000110101101000",
						 "000111000000001010100000",
						 "000111000000001101011000",
						 "000111000000010000010000",
						 "000111000000010011001000",
						 "000111000000010110000000",
						 "000111000000011000111000",
						 "000111000000011011110000",
						 "000111000000011110101000",
						 "000111000000100001100000",
						 "000111000000100100011000",
						 "000111000000100111010000",
						 "000111000000101010001000",
						 "000111000000101101000000",
						 "000111000000101111111000",
						 "000111000000110010110000",
						 "000111000000110101101000",
						 "000111000010101101011110",
						 "000111000010110000010110",
						 "000111000010110011001110",
						 "000111000010110110000110",
						 "000111000010111000111110",
						 "000111000010111011110110",
						 "000111000010111110101110",
						 "000111000011000001100110",
						 "000111000011000100011110",
						 "000111000011000111010110",
						 "000111000011001010001110",
						 "000111000011001101000110",
						 "000111000011001111111110",
						 "000111000011010010110110",
						 "000111000011010101101110",
						 "000111000011011000100110",
						 "000111000010101101011110",
						 "000111000010110000010101",
						 "000111000010110011001100",
						 "000111000010110110000011",
						 "000111000010111000111010",
						 "000111000010111011110001",
						 "000111000010111110101000",
						 "000111000011000001011111",
						 "000111000011000100010110",
						 "000111000011000111001101",
						 "000111000011001010000100",
						 "000111000011001100111011",
						 "000111000011001111110010",
						 "000111000011010010101001",
						 "000111000011010101100000",
						 "000111000011011000010111",
						 "000111000010101101011110",
						 "000111000010110000010101",
						 "000111000010110011001100",
						 "000111000010110110000011",
						 "000111000010111000111010",
						 "000111000010111011110001",
						 "000111000010111110101000",
						 "000111000011000001011111",
						 "000111000011000100010110",
						 "000111000011000111001101",
						 "000111000011001010000100",
						 "000111000011001100111011",
						 "000111000011001111110010",
						 "000111000011010010101001",
						 "000111000011010101100000",
						 "000111000011011000010111",
						 "000111000101010000011100",
						 "000111000101010011010011",
						 "000111000101010110001010",
						 "000111000101011001000001",
						 "000111000101011011111000",
						 "000111000101011110101111",
						 "000111000101100001100110",
						 "000111000101100100011101",
						 "000111000101100111010100",
						 "000111000101101010001011",
						 "000111000101101101000010",
						 "000111000101101111111001",
						 "000111000101110010110000",
						 "000111000101110101100111",
						 "000111000101111000011110",
						 "000111000101111011010101",
						 "000111000101010000011100",
						 "000111000101010011010011",
						 "000111000101010110001010",
						 "000111000101011001000001",
						 "000111000101011011111000",
						 "000111000101011110101111",
						 "000111000101100001100110",
						 "000111000101100100011101",
						 "000111000101100111010100",
						 "000111000101101010001011",
						 "000111000101101101000010",
						 "000111000101101111111001",
						 "000111000101110010110000",
						 "000111000101110101100111",
						 "000111000101111000011110",
						 "000111000101111011010101",
						 "000111000101010000011100",
						 "000111000101010011010010",
						 "000111000101010110001000",
						 "000111000101011000111110",
						 "000111000101011011110100",
						 "000111000101011110101010",
						 "000111000101100001100000",
						 "000111000101100100010110",
						 "000111000101100111001100",
						 "000111000101101010000010",
						 "000111000101101100111000",
						 "000111000101101111101110",
						 "000111000101110010100100",
						 "000111000101110101011010",
						 "000111000101111000010000",
						 "000111000101111011000110",
						 "000111000101010000011100",
						 "000111000101010011010010",
						 "000111000101010110001000",
						 "000111000101011000111110",
						 "000111000101011011110100",
						 "000111000101011110101010",
						 "000111000101100001100000",
						 "000111000101100100010110",
						 "000111000101100111001100",
						 "000111000101101010000010",
						 "000111000101101100111000",
						 "000111000101101111101110",
						 "000111000101110010100100",
						 "000111000101110101011010",
						 "000111000101111000010000",
						 "000111000101111011000110",
						 "000111000111110011011010",
						 "000111000111110110010000",
						 "000111000111111001000110",
						 "000111000111111011111100",
						 "000111000111111110110010",
						 "000111001000000001101000",
						 "000111001000000100011110",
						 "000111001000000111010100",
						 "000111001000001010001010",
						 "000111001000001101000000",
						 "000111001000001111110110",
						 "000111001000010010101100",
						 "000111001000010101100010",
						 "000111001000011000011000",
						 "000111001000011011001110",
						 "000111001000011110000100",
						 "000111000111110011011010",
						 "000111000111110110010000",
						 "000111000111111001000110",
						 "000111000111111011111100",
						 "000111000111111110110010",
						 "000111001000000001101000",
						 "000111001000000100011110",
						 "000111001000000111010100",
						 "000111001000001010001010",
						 "000111001000001101000000",
						 "000111001000001111110110",
						 "000111001000010010101100",
						 "000111001000010101100010",
						 "000111001000011000011000",
						 "000111001000011011001110",
						 "000111001000011110000100",
						 "000111000111110011011010",
						 "000111000111110110001111",
						 "000111000111111001000100",
						 "000111000111111011111001",
						 "000111000111111110101110",
						 "000111001000000001100011",
						 "000111001000000100011000",
						 "000111001000000111001101",
						 "000111001000001010000010",
						 "000111001000001100110111",
						 "000111001000001111101100",
						 "000111001000010010100001",
						 "000111001000010101010110",
						 "000111001000011000001011",
						 "000111001000011011000000",
						 "000111001000011101110101",
						 "000111000111110011011010",
						 "000111000111110110001111",
						 "000111000111111001000100",
						 "000111000111111011111001",
						 "000111000111111110101110",
						 "000111001000000001100011",
						 "000111001000000100011000",
						 "000111001000000111001101",
						 "000111001000001010000010",
						 "000111001000001100110111",
						 "000111001000001111101100",
						 "000111001000010010100001",
						 "000111001000010101010110",
						 "000111001000011000001011",
						 "000111001000011011000000",
						 "000111001000011101110101",
						 "000111001010010110011000",
						 "000111001010011001001101",
						 "000111001010011100000010",
						 "000111001010011110110111",
						 "000111001010100001101100",
						 "000111001010100100100001",
						 "000111001010100111010110",
						 "000111001010101010001011",
						 "000111001010101101000000",
						 "000111001010101111110101",
						 "000111001010110010101010",
						 "000111001010110101011111",
						 "000111001010111000010100",
						 "000111001010111011001001",
						 "000111001010111101111110",
						 "000111001011000000110011",
						 "000111001010010110011000",
						 "000111001010011001001100",
						 "000111001010011100000000",
						 "000111001010011110110100",
						 "000111001010100001101000",
						 "000111001010100100011100",
						 "000111001010100111010000",
						 "000111001010101010000100",
						 "000111001010101100111000",
						 "000111001010101111101100",
						 "000111001010110010100000",
						 "000111001010110101010100",
						 "000111001010111000001000",
						 "000111001010111010111100",
						 "000111001010111101110000",
						 "000111001011000000100100",
						 "000111001010010110011000",
						 "000111001010011001001100",
						 "000111001010011100000000",
						 "000111001010011110110100",
						 "000111001010100001101000",
						 "000111001010100100011100",
						 "000111001010100111010000",
						 "000111001010101010000100",
						 "000111001010101100111000",
						 "000111001010101111101100",
						 "000111001010110010100000",
						 "000111001010110101010100",
						 "000111001010111000001000",
						 "000111001010111010111100",
						 "000111001010111101110000",
						 "000111001011000000100100",
						 "000111001100111001010110",
						 "000111001100111100001010",
						 "000111001100111110111110",
						 "000111001101000001110010",
						 "000111001101000100100110",
						 "000111001101000111011010",
						 "000111001101001010001110",
						 "000111001101001101000010",
						 "000111001101001111110110",
						 "000111001101010010101010",
						 "000111001101010101011110",
						 "000111001101011000010010",
						 "000111001101011011000110",
						 "000111001101011101111010",
						 "000111001101100000101110",
						 "000111001101100011100010",
						 "000111001100111001010110",
						 "000111001100111100001010",
						 "000111001100111110111110",
						 "000111001101000001110010",
						 "000111001101000100100110",
						 "000111001101000111011010",
						 "000111001101001010001110",
						 "000111001101001101000010",
						 "000111001101001111110110",
						 "000111001101010010101010",
						 "000111001101010101011110",
						 "000111001101011000010010",
						 "000111001101011011000110",
						 "000111001101011101111010",
						 "000111001101100000101110",
						 "000111001101100011100010",
						 "000111001100111001010110",
						 "000111001100111100001001",
						 "000111001100111110111100",
						 "000111001101000001101111",
						 "000111001101000100100010",
						 "000111001101000111010101",
						 "000111001101001010001000",
						 "000111001101001100111011",
						 "000111001101001111101110",
						 "000111001101010010100001",
						 "000111001101010101010100",
						 "000111001101011000000111",
						 "000111001101011010111010",
						 "000111001101011101101101",
						 "000111001101100000100000",
						 "000111001101100011010011",
						 "000111001100111001010110",
						 "000111001100111100001001",
						 "000111001100111110111100",
						 "000111001101000001101111",
						 "000111001101000100100010",
						 "000111001101000111010101",
						 "000111001101001010001000",
						 "000111001101001100111011",
						 "000111001101001111101110",
						 "000111001101010010100001",
						 "000111001101010101010100",
						 "000111001101011000000111",
						 "000111001101011010111010",
						 "000111001101011101101101",
						 "000111001101100000100000",
						 "000111001101100011010011",
						 "000111001111011100010100",
						 "000111001111011111000111",
						 "000111001111100001111010",
						 "000111001111100100101101",
						 "000111001111100111100000",
						 "000111001111101010010011",
						 "000111001111101101000110",
						 "000111001111101111111001",
						 "000111001111110010101100",
						 "000111001111110101011111",
						 "000111001111111000010010",
						 "000111001111111011000101",
						 "000111001111111101111000",
						 "000111010000000000101011",
						 "000111010000000011011110",
						 "000111010000000110010001",
						 "000111001111011100010100",
						 "000111001111011111000111",
						 "000111001111100001111010",
						 "000111001111100100101101",
						 "000111001111100111100000",
						 "000111001111101010010011",
						 "000111001111101101000110",
						 "000111001111101111111001",
						 "000111001111110010101100",
						 "000111001111110101011111",
						 "000111001111111000010010",
						 "000111001111111011000101",
						 "000111001111111101111000",
						 "000111010000000000101011",
						 "000111010000000011011110",
						 "000111010000000110010001",
						 "000111001111011100010100",
						 "000111001111011111000110",
						 "000111001111100001111000",
						 "000111001111100100101010",
						 "000111001111100111011100",
						 "000111001111101010001110",
						 "000111001111101101000000",
						 "000111001111101111110010",
						 "000111001111110010100100",
						 "000111001111110101010110",
						 "000111001111111000001000",
						 "000111001111111010111010",
						 "000111001111111101101100",
						 "000111010000000000011110",
						 "000111010000000011010000",
						 "000111010000000110000010",
						 "000111010001111111010010",
						 "000111010010000010000100",
						 "000111010010000100110110",
						 "000111010010000111101000",
						 "000111010010001010011010",
						 "000111010010001101001100",
						 "000111010010001111111110",
						 "000111010010010010110000",
						 "000111010010010101100010",
						 "000111010010011000010100",
						 "000111010010011011000110",
						 "000111010010011101111000",
						 "000111010010100000101010",
						 "000111010010100011011100",
						 "000111010010100110001110",
						 "000111010010101001000000",
						 "000111010001111111010010",
						 "000111010010000010000100",
						 "000111010010000100110110",
						 "000111010010000111101000",
						 "000111010010001010011010",
						 "000111010010001101001100",
						 "000111010010001111111110",
						 "000111010010010010110000",
						 "000111010010010101100010",
						 "000111010010011000010100",
						 "000111010010011011000110",
						 "000111010010011101111000",
						 "000111010010100000101010",
						 "000111010010100011011100",
						 "000111010010100110001110",
						 "000111010010101001000000",
						 "000111010001111111010010",
						 "000111010010000010000011",
						 "000111010010000100110100",
						 "000111010010000111100101",
						 "000111010010001010010110",
						 "000111010010001101000111",
						 "000111010010001111111000",
						 "000111010010010010101001",
						 "000111010010010101011010",
						 "000111010010011000001011",
						 "000111010010011010111100",
						 "000111010010011101101101",
						 "000111010010100000011110",
						 "000111010010100011001111",
						 "000111010010100110000000",
						 "000111010010101000110001",
						 "000111010001111111010010",
						 "000111010010000010000011",
						 "000111010010000100110100",
						 "000111010010000111100101",
						 "000111010010001010010110",
						 "000111010010001101000111",
						 "000111010010001111111000",
						 "000111010010010010101001",
						 "000111010010010101011010",
						 "000111010010011000001011",
						 "000111010010011010111100",
						 "000111010010011101101101",
						 "000111010010100000011110",
						 "000111010010100011001111",
						 "000111010010100110000000",
						 "000111010010101000110001",
						 "000111010100100010010000",
						 "000111010100100101000001",
						 "000111010100100111110010",
						 "000111010100101010100011",
						 "000111010100101101010100",
						 "000111010100110000000101",
						 "000111010100110010110110",
						 "000111010100110101100111",
						 "000111010100111000011000",
						 "000111010100111011001001",
						 "000111010100111101111010",
						 "000111010101000000101011",
						 "000111010101000011011100",
						 "000111010101000110001101",
						 "000111010101001000111110",
						 "000111010101001011101111",
						 "000111010100100010010000",
						 "000111010100100101000001",
						 "000111010100100111110010",
						 "000111010100101010100011",
						 "000111010100101101010100",
						 "000111010100110000000101",
						 "000111010100110010110110",
						 "000111010100110101100111",
						 "000111010100111000011000",
						 "000111010100111011001001",
						 "000111010100111101111010",
						 "000111010101000000101011",
						 "000111010101000011011100",
						 "000111010101000110001101",
						 "000111010101001000111110",
						 "000111010101001011101111",
						 "000111010100100010010000",
						 "000111010100100101000000",
						 "000111010100100111110000",
						 "000111010100101010100000",
						 "000111010100101101010000",
						 "000111010100110000000000",
						 "000111010100110010110000",
						 "000111010100110101100000",
						 "000111010100111000010000",
						 "000111010100111011000000",
						 "000111010100111101110000",
						 "000111010101000000100000",
						 "000111010101000011010000",
						 "000111010101000110000000",
						 "000111010101001000110000",
						 "000111010101001011100000",
						 "000111010100100010010000",
						 "000111010100100101000000",
						 "000111010100100111110000",
						 "000111010100101010100000",
						 "000111010100101101010000",
						 "000111010100110000000000",
						 "000111010100110010110000",
						 "000111010100110101100000",
						 "000111010100111000010000",
						 "000111010100111011000000",
						 "000111010100111101110000",
						 "000111010101000000100000",
						 "000111010101000011010000",
						 "000111010101000110000000",
						 "000111010101001000110000",
						 "000111010101001011100000",
						 "000111010111000101001110",
						 "000111010111000111111110",
						 "000111010111001010101110",
						 "000111010111001101011110",
						 "000111010111010000001110",
						 "000111010111010010111110",
						 "000111010111010101101110",
						 "000111010111011000011110",
						 "000111010111011011001110",
						 "000111010111011101111110",
						 "000111010111100000101110",
						 "000111010111100011011110",
						 "000111010111100110001110",
						 "000111010111101000111110",
						 "000111010111101011101110",
						 "000111010111101110011110",
						 "000111010111000101001110",
						 "000111010111000111111101",
						 "000111010111001010101100",
						 "000111010111001101011011",
						 "000111010111010000001010",
						 "000111010111010010111001",
						 "000111010111010101101000",
						 "000111010111011000010111",
						 "000111010111011011000110",
						 "000111010111011101110101",
						 "000111010111100000100100",
						 "000111010111100011010011",
						 "000111010111100110000010",
						 "000111010111101000110001",
						 "000111010111101011100000",
						 "000111010111101110001111",
						 "000111010111000101001110",
						 "000111010111000111111101",
						 "000111010111001010101100",
						 "000111010111001101011011",
						 "000111010111010000001010",
						 "000111010111010010111001",
						 "000111010111010101101000",
						 "000111010111011000010111",
						 "000111010111011011000110",
						 "000111010111011101110101",
						 "000111010111100000100100",
						 "000111010111100011010011",
						 "000111010111100110000010",
						 "000111010111101000110001",
						 "000111010111101011100000",
						 "000111010111101110001111",
						 "000111010111000101001110",
						 "000111010111000111111101",
						 "000111010111001010101100",
						 "000111010111001101011011",
						 "000111010111010000001010",
						 "000111010111010010111001",
						 "000111010111010101101000",
						 "000111010111011000010111",
						 "000111010111011011000110",
						 "000111010111011101110101",
						 "000111010111100000100100",
						 "000111010111100011010011",
						 "000111010111100110000010",
						 "000111010111101000110001",
						 "000111010111101011100000",
						 "000111010111101110001111",
						 "000111011001101000001100",
						 "000111011001101010111011",
						 "000111011001101101101010",
						 "000111011001110000011001",
						 "000111011001110011001000",
						 "000111011001110101110111",
						 "000111011001111000100110",
						 "000111011001111011010101",
						 "000111011001111110000100",
						 "000111011010000000110011",
						 "000111011010000011100010",
						 "000111011010000110010001",
						 "000111011010001001000000",
						 "000111011010001011101111",
						 "000111011010001110011110",
						 "000111011010010001001101",
						 "000111011001101000001100",
						 "000111011001101010111010",
						 "000111011001101101101000",
						 "000111011001110000010110",
						 "000111011001110011000100",
						 "000111011001110101110010",
						 "000111011001111000100000",
						 "000111011001111011001110",
						 "000111011001111101111100",
						 "000111011010000000101010",
						 "000111011010000011011000",
						 "000111011010000110000110",
						 "000111011010001000110100",
						 "000111011010001011100010",
						 "000111011010001110010000",
						 "000111011010010000111110",
						 "000111011001101000001100",
						 "000111011001101010111010",
						 "000111011001101101101000",
						 "000111011001110000010110",
						 "000111011001110011000100",
						 "000111011001110101110010",
						 "000111011001111000100000",
						 "000111011001111011001110",
						 "000111011001111101111100",
						 "000111011010000000101010",
						 "000111011010000011011000",
						 "000111011010000110000110",
						 "000111011010001000110100",
						 "000111011010001011100010",
						 "000111011010001110010000",
						 "000111011010010000111110",
						 "000111011100001011001010",
						 "000111011100001101111000",
						 "000111011100010000100110",
						 "000111011100010011010100",
						 "000111011100010110000010",
						 "000111011100011000110000",
						 "000111011100011011011110",
						 "000111011100011110001100",
						 "000111011100100000111010",
						 "000111011100100011101000",
						 "000111011100100110010110",
						 "000111011100101001000100",
						 "000111011100101011110010",
						 "000111011100101110100000",
						 "000111011100110001001110",
						 "000111011100110011111100",
						 "000111011100001011001010",
						 "000111011100001101110111",
						 "000111011100010000100100",
						 "000111011100010011010001",
						 "000111011100010101111110",
						 "000111011100011000101011",
						 "000111011100011011011000",
						 "000111011100011110000101",
						 "000111011100100000110010",
						 "000111011100100011011111",
						 "000111011100100110001100",
						 "000111011100101000111001",
						 "000111011100101011100110",
						 "000111011100101110010011",
						 "000111011100110001000000",
						 "000111011100110011101101",
						 "000111011100001011001010",
						 "000111011100001101110111",
						 "000111011100010000100100",
						 "000111011100010011010001",
						 "000111011100010101111110",
						 "000111011100011000101011",
						 "000111011100011011011000",
						 "000111011100011110000101",
						 "000111011100100000110010",
						 "000111011100100011011111",
						 "000111011100100110001100",
						 "000111011100101000111001",
						 "000111011100101011100110",
						 "000111011100101110010011",
						 "000111011100110001000000",
						 "000111011100110011101101",
						 "000111011100001011001010",
						 "000111011100001101110111",
						 "000111011100010000100100",
						 "000111011100010011010001",
						 "000111011100010101111110",
						 "000111011100011000101011",
						 "000111011100011011011000",
						 "000111011100011110000101",
						 "000111011100100000110010",
						 "000111011100100011011111",
						 "000111011100100110001100",
						 "000111011100101000111001",
						 "000111011100101011100110",
						 "000111011100101110010011",
						 "000111011100110001000000",
						 "000111011100110011101101",
						 "000111011110101110001000",
						 "000111011110110000110101",
						 "000111011110110011100010",
						 "000111011110110110001111",
						 "000111011110111000111100",
						 "000111011110111011101001",
						 "000111011110111110010110",
						 "000111011111000001000011",
						 "000111011111000011110000",
						 "000111011111000110011101",
						 "000111011111001001001010",
						 "000111011111001011110111",
						 "000111011111001110100100",
						 "000111011111010001010001",
						 "000111011111010011111110",
						 "000111011111010110101011",
						 "000111011110101110001000",
						 "000111011110110000110100",
						 "000111011110110011100000",
						 "000111011110110110001100",
						 "000111011110111000111000",
						 "000111011110111011100100",
						 "000111011110111110010000",
						 "000111011111000000111100",
						 "000111011111000011101000",
						 "000111011111000110010100",
						 "000111011111001001000000",
						 "000111011111001011101100",
						 "000111011111001110011000",
						 "000111011111010001000100",
						 "000111011111010011110000",
						 "000111011111010110011100",
						 "000111011110101110001000",
						 "000111011110110000110100",
						 "000111011110110011100000",
						 "000111011110110110001100",
						 "000111011110111000111000",
						 "000111011110111011100100",
						 "000111011110111110010000",
						 "000111011111000000111100",
						 "000111011111000011101000",
						 "000111011111000110010100",
						 "000111011111001001000000",
						 "000111011111001011101100",
						 "000111011111001110011000",
						 "000111011111010001000100",
						 "000111011111010011110000",
						 "000111011111010110011100",
						 "000111011110101110001000",
						 "000111011110110000110100",
						 "000111011110110011100000",
						 "000111011110110110001100",
						 "000111011110111000111000",
						 "000111011110111011100100",
						 "000111011110111110010000",
						 "000111011111000000111100",
						 "000111011111000011101000",
						 "000111011111000110010100",
						 "000111011111001001000000",
						 "000111011111001011101100",
						 "000111011111001110011000",
						 "000111011111010001000100",
						 "000111011111010011110000",
						 "000111011111010110011100",
						 "000111100001010001000110",
						 "000111100001010011110001",
						 "000111100001010110011100",
						 "000111100001011001000111",
						 "000111100001011011110010",
						 "000111100001011110011101",
						 "000111100001100001001000",
						 "000111100001100011110011",
						 "000111100001100110011110",
						 "000111100001101001001001",
						 "000111100001101011110100",
						 "000111100001101110011111",
						 "000111100001110001001010",
						 "000111100001110011110101",
						 "000111100001110110100000",
						 "000111100001111001001011",
						 "000111100001010001000110",
						 "000111100001010011110001",
						 "000111100001010110011100",
						 "000111100001011001000111",
						 "000111100001011011110010",
						 "000111100001011110011101",
						 "000111100001100001001000",
						 "000111100001100011110011",
						 "000111100001100110011110",
						 "000111100001101001001001",
						 "000111100001101011110100",
						 "000111100001101110011111",
						 "000111100001110001001010",
						 "000111100001110011110101",
						 "000111100001110110100000",
						 "000111100001111001001011",
						 "000111100001010001000110",
						 "000111100001010011110001",
						 "000111100001010110011100",
						 "000111100001011001000111",
						 "000111100001011011110010",
						 "000111100001011110011101",
						 "000111100001100001001000",
						 "000111100001100011110011",
						 "000111100001100110011110",
						 "000111100001101001001001",
						 "000111100001101011110100",
						 "000111100001101110011111",
						 "000111100001110001001010",
						 "000111100001110011110101",
						 "000111100001110110100000",
						 "000111100001111001001011",
						 "000111100001010001000110",
						 "000111100001010011110001",
						 "000111100001010110011100",
						 "000111100001011001000111",
						 "000111100001011011110010",
						 "000111100001011110011101",
						 "000111100001100001001000",
						 "000111100001100011110011",
						 "000111100001100110011110",
						 "000111100001101001001001",
						 "000111100001101011110100",
						 "000111100001101110011111",
						 "000111100001110001001010",
						 "000111100001110011110101",
						 "000111100001110110100000",
						 "000111100001111001001011",
						 "000111100011110100000100",
						 "000111100011110110101110",
						 "000111100011111001011000",
						 "000111100011111100000010",
						 "000111100011111110101100",
						 "000111100100000001010110",
						 "000111100100000100000000",
						 "000111100100000110101010",
						 "000111100100001001010100",
						 "000111100100001011111110",
						 "000111100100001110101000",
						 "000111100100010001010010",
						 "000111100100010011111100",
						 "000111100100010110100110",
						 "000111100100011001010000",
						 "000111100100011011111010",
						 "000111100011110100000100",
						 "000111100011110110101110",
						 "000111100011111001011000",
						 "000111100011111100000010",
						 "000111100011111110101100",
						 "000111100100000001010110",
						 "000111100100000100000000",
						 "000111100100000110101010",
						 "000111100100001001010100",
						 "000111100100001011111110",
						 "000111100100001110101000",
						 "000111100100010001010010",
						 "000111100100010011111100",
						 "000111100100010110100110",
						 "000111100100011001010000",
						 "000111100100011011111010",
						 "000111100011110100000100",
						 "000111100011110110101110",
						 "000111100011111001011000",
						 "000111100011111100000010",
						 "000111100011111110101100",
						 "000111100100000001010110",
						 "000111100100000100000000",
						 "000111100100000110101010",
						 "000111100100001001010100",
						 "000111100100001011111110",
						 "000111100100001110101000",
						 "000111100100010001010010",
						 "000111100100010011111100",
						 "000111100100010110100110",
						 "000111100100011001010000",
						 "000111100100011011111010",
						 "000111100110010111000010",
						 "000111100110011001101011",
						 "000111100110011100010100",
						 "000111100110011110111101",
						 "000111100110100001100110",
						 "000111100110100100001111",
						 "000111100110100110111000",
						 "000111100110101001100001",
						 "000111100110101100001010",
						 "000111100110101110110011",
						 "000111100110110001011100",
						 "000111100110110100000101",
						 "000111100110110110101110",
						 "000111100110111001010111",
						 "000111100110111100000000",
						 "000111100110111110101001",
						 "000111100110010111000010",
						 "000111100110011001101011",
						 "000111100110011100010100",
						 "000111100110011110111101",
						 "000111100110100001100110",
						 "000111100110100100001111",
						 "000111100110100110111000",
						 "000111100110101001100001",
						 "000111100110101100001010",
						 "000111100110101110110011",
						 "000111100110110001011100",
						 "000111100110110100000101",
						 "000111100110110110101110",
						 "000111100110111001010111",
						 "000111100110111100000000",
						 "000111100110111110101001",
						 "000111100110010111000010",
						 "000111100110011001101011",
						 "000111100110011100010100",
						 "000111100110011110111101",
						 "000111100110100001100110",
						 "000111100110100100001111",
						 "000111100110100110111000",
						 "000111100110101001100001",
						 "000111100110101100001010",
						 "000111100110101110110011",
						 "000111100110110001011100",
						 "000111100110110100000101",
						 "000111100110110110101110",
						 "000111100110111001010111",
						 "000111100110111100000000",
						 "000111100110111110101001",
						 "000111100110010111000010",
						 "000111100110011001101010",
						 "000111100110011100010010",
						 "000111100110011110111010",
						 "000111100110100001100010",
						 "000111100110100100001010",
						 "000111100110100110110010",
						 "000111100110101001011010",
						 "000111100110101100000010",
						 "000111100110101110101010",
						 "000111100110110001010010",
						 "000111100110110011111010",
						 "000111100110110110100010",
						 "000111100110111001001010",
						 "000111100110111011110010",
						 "000111100110111110011010",
						 "000111101000111010000000",
						 "000111101000111100101000",
						 "000111101000111111010000",
						 "000111101001000001111000",
						 "000111101001000100100000",
						 "000111101001000111001000",
						 "000111101001001001110000",
						 "000111101001001100011000",
						 "000111101001001111000000",
						 "000111101001010001101000",
						 "000111101001010100010000",
						 "000111101001010110111000",
						 "000111101001011001100000",
						 "000111101001011100001000",
						 "000111101001011110110000",
						 "000111101001100001011000",
						 "000111101000111010000000",
						 "000111101000111100101000",
						 "000111101000111111010000",
						 "000111101001000001111000",
						 "000111101001000100100000",
						 "000111101001000111001000",
						 "000111101001001001110000",
						 "000111101001001100011000",
						 "000111101001001111000000",
						 "000111101001010001101000",
						 "000111101001010100010000",
						 "000111101001010110111000",
						 "000111101001011001100000",
						 "000111101001011100001000",
						 "000111101001011110110000",
						 "000111101001100001011000",
						 "000111101000111010000000",
						 "000111101000111100101000",
						 "000111101000111111010000",
						 "000111101001000001111000",
						 "000111101001000100100000",
						 "000111101001000111001000",
						 "000111101001001001110000",
						 "000111101001001100011000",
						 "000111101001001111000000",
						 "000111101001010001101000",
						 "000111101001010100010000",
						 "000111101001010110111000",
						 "000111101001011001100000",
						 "000111101001011100001000",
						 "000111101001011110110000",
						 "000111101001100001011000",
						 "000111101000111010000000",
						 "000111101000111100100111",
						 "000111101000111111001110",
						 "000111101001000001110101",
						 "000111101001000100011100",
						 "000111101001000111000011",
						 "000111101001001001101010",
						 "000111101001001100010001",
						 "000111101001001110111000",
						 "000111101001010001011111",
						 "000111101001010100000110",
						 "000111101001010110101101",
						 "000111101001011001010100",
						 "000111101001011011111011",
						 "000111101001011110100010",
						 "000111101001100001001001",
						 "000111101011011100111110",
						 "000111101011011111100101",
						 "000111101011100010001100",
						 "000111101011100100110011",
						 "000111101011100111011010",
						 "000111101011101010000001",
						 "000111101011101100101000",
						 "000111101011101111001111",
						 "000111101011110001110110",
						 "000111101011110100011101",
						 "000111101011110111000100",
						 "000111101011111001101011",
						 "000111101011111100010010",
						 "000111101011111110111001",
						 "000111101100000001100000",
						 "000111101100000100000111",
						 "000111101011011100111110",
						 "000111101011011111100101",
						 "000111101011100010001100",
						 "000111101011100100110011",
						 "000111101011100111011010",
						 "000111101011101010000001",
						 "000111101011101100101000",
						 "000111101011101111001111",
						 "000111101011110001110110",
						 "000111101011110100011101",
						 "000111101011110111000100",
						 "000111101011111001101011",
						 "000111101011111100010010",
						 "000111101011111110111001",
						 "000111101100000001100000",
						 "000111101100000100000111",
						 "000111101011011100111110",
						 "000111101011011111100100",
						 "000111101011100010001010",
						 "000111101011100100110000",
						 "000111101011100111010110",
						 "000111101011101001111100",
						 "000111101011101100100010",
						 "000111101011101111001000",
						 "000111101011110001101110",
						 "000111101011110100010100",
						 "000111101011110110111010",
						 "000111101011111001100000",
						 "000111101011111100000110",
						 "000111101011111110101100",
						 "000111101100000001010010",
						 "000111101100000011111000",
						 "000111101011011100111110",
						 "000111101011011111100100",
						 "000111101011100010001010",
						 "000111101011100100110000",
						 "000111101011100111010110",
						 "000111101011101001111100",
						 "000111101011101100100010",
						 "000111101011101111001000",
						 "000111101011110001101110",
						 "000111101011110100010100",
						 "000111101011110110111010",
						 "000111101011111001100000",
						 "000111101011111100000110",
						 "000111101011111110101100",
						 "000111101100000001010010",
						 "000111101100000011111000",
						 "000111101101111111111100",
						 "000111101110000010100010",
						 "000111101110000101001000",
						 "000111101110000111101110",
						 "000111101110001010010100",
						 "000111101110001100111010",
						 "000111101110001111100000",
						 "000111101110010010000110",
						 "000111101110010100101100",
						 "000111101110010111010010",
						 "000111101110011001111000",
						 "000111101110011100011110",
						 "000111101110011111000100",
						 "000111101110100001101010",
						 "000111101110100100010000",
						 "000111101110100110110110",
						 "000111101101111111111100",
						 "000111101110000010100010",
						 "000111101110000101001000",
						 "000111101110000111101110",
						 "000111101110001010010100",
						 "000111101110001100111010",
						 "000111101110001111100000",
						 "000111101110010010000110",
						 "000111101110010100101100",
						 "000111101110010111010010",
						 "000111101110011001111000",
						 "000111101110011100011110",
						 "000111101110011111000100",
						 "000111101110100001101010",
						 "000111101110100100010000",
						 "000111101110100110110110",
						 "000111101101111111111100",
						 "000111101110000010100001",
						 "000111101110000101000110",
						 "000111101110000111101011",
						 "000111101110001010010000",
						 "000111101110001100110101",
						 "000111101110001111011010",
						 "000111101110010001111111",
						 "000111101110010100100100",
						 "000111101110010111001001",
						 "000111101110011001101110",
						 "000111101110011100010011",
						 "000111101110011110111000",
						 "000111101110100001011101",
						 "000111101110100100000010",
						 "000111101110100110100111",
						 "000111101101111111111100",
						 "000111101110000010100001",
						 "000111101110000101000110",
						 "000111101110000111101011",
						 "000111101110001010010000",
						 "000111101110001100110101",
						 "000111101110001111011010",
						 "000111101110010001111111",
						 "000111101110010100100100",
						 "000111101110010111001001",
						 "000111101110011001101110",
						 "000111101110011100010011",
						 "000111101110011110111000",
						 "000111101110100001011101",
						 "000111101110100100000010",
						 "000111101110100110100111",
						 "000111110000100010111010",
						 "000111110000100101011111",
						 "000111110000101000000100",
						 "000111110000101010101001",
						 "000111110000101101001110",
						 "000111110000101111110011",
						 "000111110000110010011000",
						 "000111110000110100111101",
						 "000111110000110111100010",
						 "000111110000111010000111",
						 "000111110000111100101100",
						 "000111110000111111010001",
						 "000111110001000001110110",
						 "000111110001000100011011",
						 "000111110001000111000000",
						 "000111110001001001100101",
						 "000111110000100010111010",
						 "000111110000100101011110",
						 "000111110000101000000010",
						 "000111110000101010100110",
						 "000111110000101101001010",
						 "000111110000101111101110",
						 "000111110000110010010010",
						 "000111110000110100110110",
						 "000111110000110111011010",
						 "000111110000111001111110",
						 "000111110000111100100010",
						 "000111110000111111000110",
						 "000111110001000001101010",
						 "000111110001000100001110",
						 "000111110001000110110010",
						 "000111110001001001010110",
						 "000111110000100010111010",
						 "000111110000100101011110",
						 "000111110000101000000010",
						 "000111110000101010100110",
						 "000111110000101101001010",
						 "000111110000101111101110",
						 "000111110000110010010010",
						 "000111110000110100110110",
						 "000111110000110111011010",
						 "000111110000111001111110",
						 "000111110000111100100010",
						 "000111110000111111000110",
						 "000111110001000001101010",
						 "000111110001000100001110",
						 "000111110001000110110010",
						 "000111110001001001010110",
						 "000111110000100010111010",
						 "000111110000100101011110",
						 "000111110000101000000010",
						 "000111110000101010100110",
						 "000111110000101101001010",
						 "000111110000101111101110",
						 "000111110000110010010010",
						 "000111110000110100110110",
						 "000111110000110111011010",
						 "000111110000111001111110",
						 "000111110000111100100010",
						 "000111110000111111000110",
						 "000111110001000001101010",
						 "000111110001000100001110",
						 "000111110001000110110010",
						 "000111110001001001010110",
						 "000111110011000101111000",
						 "000111110011001000011011",
						 "000111110011001010111110",
						 "000111110011001101100001",
						 "000111110011010000000100",
						 "000111110011010010100111",
						 "000111110011010101001010",
						 "000111110011010111101101",
						 "000111110011011010010000",
						 "000111110011011100110011",
						 "000111110011011111010110",
						 "000111110011100001111001",
						 "000111110011100100011100",
						 "000111110011100110111111",
						 "000111110011101001100010",
						 "000111110011101100000101",
						 "000111110011000101111000",
						 "000111110011001000011011",
						 "000111110011001010111110",
						 "000111110011001101100001",
						 "000111110011010000000100",
						 "000111110011010010100111",
						 "000111110011010101001010",
						 "000111110011010111101101",
						 "000111110011011010010000",
						 "000111110011011100110011",
						 "000111110011011111010110",
						 "000111110011100001111001",
						 "000111110011100100011100",
						 "000111110011100110111111",
						 "000111110011101001100010",
						 "000111110011101100000101",
						 "000111110011000101111000",
						 "000111110011001000011011",
						 "000111110011001010111110",
						 "000111110011001101100001",
						 "000111110011010000000100",
						 "000111110011010010100111",
						 "000111110011010101001010",
						 "000111110011010111101101",
						 "000111110011011010010000",
						 "000111110011011100110011",
						 "000111110011011111010110",
						 "000111110011100001111001",
						 "000111110011100100011100",
						 "000111110011100110111111",
						 "000111110011101001100010",
						 "000111110011101100000101",
						 "000111110011000101111000",
						 "000111110011001000011011",
						 "000111110011001010111110",
						 "000111110011001101100001",
						 "000111110011010000000100",
						 "000111110011010010100111",
						 "000111110011010101001010",
						 "000111110011010111101101",
						 "000111110011011010010000",
						 "000111110011011100110011",
						 "000111110011011111010110",
						 "000111110011100001111001",
						 "000111110011100100011100",
						 "000111110011100110111111",
						 "000111110011101001100010",
						 "000111110011101100000101",
						 "000111110101101000110110",
						 "000111110101101011011000",
						 "000111110101101101111010",
						 "000111110101110000011100",
						 "000111110101110010111110",
						 "000111110101110101100000",
						 "000111110101111000000010",
						 "000111110101111010100100",
						 "000111110101111101000110",
						 "000111110101111111101000",
						 "000111110110000010001010",
						 "000111110110000100101100",
						 "000111110110000111001110",
						 "000111110110001001110000",
						 "000111110110001100010010",
						 "000111110110001110110100",
						 "000111110101101000110110",
						 "000111110101101011011000",
						 "000111110101101101111010",
						 "000111110101110000011100",
						 "000111110101110010111110",
						 "000111110101110101100000",
						 "000111110101111000000010",
						 "000111110101111010100100",
						 "000111110101111101000110",
						 "000111110101111111101000",
						 "000111110110000010001010",
						 "000111110110000100101100",
						 "000111110110000111001110",
						 "000111110110001001110000",
						 "000111110110001100010010",
						 "000111110110001110110100",
						 "000111110101101000110110",
						 "000111110101101011011000",
						 "000111110101101101111010",
						 "000111110101110000011100",
						 "000111110101110010111110",
						 "000111110101110101100000",
						 "000111110101111000000010",
						 "000111110101111010100100",
						 "000111110101111101000110",
						 "000111110101111111101000",
						 "000111110110000010001010",
						 "000111110110000100101100",
						 "000111110110000111001110",
						 "000111110110001001110000",
						 "000111110110001100010010",
						 "000111110110001110110100",
						 "000111110101101000110110",
						 "000111110101101011010111",
						 "000111110101101101111000",
						 "000111110101110000011001",
						 "000111110101110010111010",
						 "000111110101110101011011",
						 "000111110101110111111100",
						 "000111110101111010011101",
						 "000111110101111100111110",
						 "000111110101111111011111",
						 "000111110110000010000000",
						 "000111110110000100100001",
						 "000111110110000111000010",
						 "000111110110001001100011",
						 "000111110110001100000100",
						 "000111110110001110100101",
						 "000111111000001011110100",
						 "000111111000001110010101",
						 "000111111000010000110110",
						 "000111111000010011010111",
						 "000111111000010101111000",
						 "000111111000011000011001",
						 "000111111000011010111010",
						 "000111111000011101011011",
						 "000111111000011111111100",
						 "000111111000100010011101",
						 "000111111000100100111110",
						 "000111111000100111011111",
						 "000111111000101010000000",
						 "000111111000101100100001",
						 "000111111000101111000010",
						 "000111111000110001100011",
						 "000111111000001011110100",
						 "000111111000001110010101",
						 "000111111000010000110110",
						 "000111111000010011010111",
						 "000111111000010101111000",
						 "000111111000011000011001",
						 "000111111000011010111010",
						 "000111111000011101011011",
						 "000111111000011111111100",
						 "000111111000100010011101",
						 "000111111000100100111110",
						 "000111111000100111011111",
						 "000111111000101010000000",
						 "000111111000101100100001",
						 "000111111000101111000010",
						 "000111111000110001100011",
						 "000111111000001011110100",
						 "000111111000001110010100",
						 "000111111000010000110100",
						 "000111111000010011010100",
						 "000111111000010101110100",
						 "000111111000011000010100",
						 "000111111000011010110100",
						 "000111111000011101010100",
						 "000111111000011111110100",
						 "000111111000100010010100",
						 "000111111000100100110100",
						 "000111111000100111010100",
						 "000111111000101001110100",
						 "000111111000101100010100",
						 "000111111000101110110100",
						 "000111111000110001010100",
						 "000111111000001011110100",
						 "000111111000001110010100",
						 "000111111000010000110100",
						 "000111111000010011010100",
						 "000111111000010101110100",
						 "000111111000011000010100",
						 "000111111000011010110100",
						 "000111111000011101010100",
						 "000111111000011111110100",
						 "000111111000100010010100",
						 "000111111000100100110100",
						 "000111111000100111010100",
						 "000111111000101001110100",
						 "000111111000101100010100",
						 "000111111000101110110100",
						 "000111111000110001010100",
						 "000111111010101110110010",
						 "000111111010110001010010",
						 "000111111010110011110010",
						 "000111111010110110010010",
						 "000111111010111000110010",
						 "000111111010111011010010",
						 "000111111010111101110010",
						 "000111111011000000010010",
						 "000111111011000010110010",
						 "000111111011000101010010",
						 "000111111011000111110010",
						 "000111111011001010010010",
						 "000111111011001100110010",
						 "000111111011001111010010",
						 "000111111011010001110010",
						 "000111111011010100010010",
						 "000111111010101110110010",
						 "000111111010110001010001",
						 "000111111010110011110000",
						 "000111111010110110001111",
						 "000111111010111000101110",
						 "000111111010111011001101",
						 "000111111010111101101100",
						 "000111111011000000001011",
						 "000111111011000010101010",
						 "000111111011000101001001",
						 "000111111011000111101000",
						 "000111111011001010000111",
						 "000111111011001100100110",
						 "000111111011001111000101",
						 "000111111011010001100100",
						 "000111111011010100000011",
						 "000111111010101110110010",
						 "000111111010110001010001",
						 "000111111010110011110000",
						 "000111111010110110001111",
						 "000111111010111000101110",
						 "000111111010111011001101",
						 "000111111010111101101100",
						 "000111111011000000001011",
						 "000111111011000010101010",
						 "000111111011000101001001",
						 "000111111011000111101000",
						 "000111111011001010000111",
						 "000111111011001100100110",
						 "000111111011001111000101",
						 "000111111011010001100100",
						 "000111111011010100000011",
						 "000111111010101110110010",
						 "000111111010110001010001",
						 "000111111010110011110000",
						 "000111111010110110001111",
						 "000111111010111000101110",
						 "000111111010111011001101",
						 "000111111010111101101100",
						 "000111111011000000001011",
						 "000111111011000010101010",
						 "000111111011000101001001",
						 "000111111011000111101000",
						 "000111111011001010000111",
						 "000111111011001100100110",
						 "000111111011001111000101",
						 "000111111011010001100100",
						 "000111111011010100000011",
						 "000111111101010001110000",
						 "000111111101010100001111",
						 "000111111101010110101110",
						 "000111111101011001001101",
						 "000111111101011011101100",
						 "000111111101011110001011",
						 "000111111101100000101010",
						 "000111111101100011001001",
						 "000111111101100101101000",
						 "000111111101101000000111",
						 "000111111101101010100110",
						 "000111111101101101000101",
						 "000111111101101111100100",
						 "000111111101110010000011",
						 "000111111101110100100010",
						 "000111111101110111000001",
						 "000111111101010001110000",
						 "000111111101010100001110",
						 "000111111101010110101100",
						 "000111111101011001001010",
						 "000111111101011011101000",
						 "000111111101011110000110",
						 "000111111101100000100100",
						 "000111111101100011000010",
						 "000111111101100101100000",
						 "000111111101100111111110",
						 "000111111101101010011100",
						 "000111111101101100111010",
						 "000111111101101111011000",
						 "000111111101110001110110",
						 "000111111101110100010100",
						 "000111111101110110110010",
						 "000111111101010001110000",
						 "000111111101010100001110",
						 "000111111101010110101100",
						 "000111111101011001001010",
						 "000111111101011011101000",
						 "000111111101011110000110",
						 "000111111101100000100100",
						 "000111111101100011000010",
						 "000111111101100101100000",
						 "000111111101100111111110",
						 "000111111101101010011100",
						 "000111111101101100111010",
						 "000111111101101111011000",
						 "000111111101110001110110",
						 "000111111101110100010100",
						 "000111111101110110110010",
						 "000111111101010001110000",
						 "000111111101010100001110",
						 "000111111101010110101100",
						 "000111111101011001001010",
						 "000111111101011011101000",
						 "000111111101011110000110",
						 "000111111101100000100100",
						 "000111111101100011000010",
						 "000111111101100101100000",
						 "000111111101100111111110",
						 "000111111101101010011100",
						 "000111111101101100111010",
						 "000111111101101111011000",
						 "000111111101110001110110",
						 "000111111101110100010100",
						 "000111111101110110110010",
						 "000111111111110100101110",
						 "000111111111110111001011",
						 "000111111111111001101000",
						 "000111111111111100000101",
						 "000111111111111110100010",
						 "001000000000000000111111",
						 "001000000000000011011100",
						 "001000000000000101111001",
						 "001000000000001000010110",
						 "001000000000001010110011",
						 "001000000000001101010000",
						 "001000000000001111101101",
						 "001000000000010010001010",
						 "001000000000010100100111",
						 "001000000000010111000100",
						 "001000000000011001100001",
						 "000111111111110100101110",
						 "000111111111110111001011",
						 "000111111111111001101000",
						 "000111111111111100000101",
						 "000111111111111110100010",
						 "001000000000000000111111",
						 "001000000000000011011100",
						 "001000000000000101111001",
						 "001000000000001000010110",
						 "001000000000001010110011",
						 "001000000000001101010000",
						 "001000000000001111101101",
						 "001000000000010010001010",
						 "001000000000010100100111",
						 "001000000000010111000100",
						 "001000000000011001100001",
						 "000111111111110100101110",
						 "000111111111110111001011",
						 "000111111111111001101000",
						 "000111111111111100000101",
						 "000111111111111110100010",
						 "001000000000000000111111",
						 "001000000000000011011100",
						 "001000000000000101111001",
						 "001000000000001000010110",
						 "001000000000001010110011",
						 "001000000000001101010000",
						 "001000000000001111101101",
						 "001000000000010010001010",
						 "001000000000010100100111",
						 "001000000000010111000100",
						 "001000000000011001100001",
						 "000111111111110100101110",
						 "000111111111110111001010",
						 "000111111111111001100110",
						 "000111111111111100000010",
						 "000111111111111110011110",
						 "001000000000000000111010",
						 "001000000000000011010110",
						 "001000000000000101110010",
						 "001000000000001000001110",
						 "001000000000001010101010",
						 "001000000000001101000110",
						 "001000000000001111100010",
						 "001000000000010001111110",
						 "001000000000010100011010",
						 "001000000000010110110110",
						 "001000000000011001010010",
						 "001000000010010111101100",
						 "001000000010011010001000",
						 "001000000010011100100100",
						 "001000000010011111000000",
						 "001000000010100001011100",
						 "001000000010100011111000",
						 "001000000010100110010100",
						 "001000000010101000110000",
						 "001000000010101011001100",
						 "001000000010101101101000",
						 "001000000010110000000100",
						 "001000000010110010100000",
						 "001000000010110100111100",
						 "001000000010110111011000",
						 "001000000010111001110100",
						 "001000000010111100010000",
						 "001000000010010111101100",
						 "001000000010011010001000",
						 "001000000010011100100100",
						 "001000000010011111000000",
						 "001000000010100001011100",
						 "001000000010100011111000",
						 "001000000010100110010100",
						 "001000000010101000110000",
						 "001000000010101011001100",
						 "001000000010101101101000",
						 "001000000010110000000100",
						 "001000000010110010100000",
						 "001000000010110100111100",
						 "001000000010110111011000",
						 "001000000010111001110100",
						 "001000000010111100010000",
						 "001000000010010111101100",
						 "001000000010011010000111",
						 "001000000010011100100010",
						 "001000000010011110111101",
						 "001000000010100001011000",
						 "001000000010100011110011",
						 "001000000010100110001110",
						 "001000000010101000101001",
						 "001000000010101011000100",
						 "001000000010101101011111",
						 "001000000010101111111010",
						 "001000000010110010010101",
						 "001000000010110100110000",
						 "001000000010110111001011",
						 "001000000010111001100110",
						 "001000000010111100000001",
						 "001000000010010111101100",
						 "001000000010011010000111",
						 "001000000010011100100010",
						 "001000000010011110111101",
						 "001000000010100001011000",
						 "001000000010100011110011",
						 "001000000010100110001110",
						 "001000000010101000101001",
						 "001000000010101011000100",
						 "001000000010101101011111",
						 "001000000010101111111010",
						 "001000000010110010010101",
						 "001000000010110100110000",
						 "001000000010110111001011",
						 "001000000010111001100110",
						 "001000000010111100000001",
						 "001000000010010111101100",
						 "001000000010011010000111",
						 "001000000010011100100010",
						 "001000000010011110111101",
						 "001000000010100001011000",
						 "001000000010100011110011",
						 "001000000010100110001110",
						 "001000000010101000101001",
						 "001000000010101011000100",
						 "001000000010101101011111",
						 "001000000010101111111010",
						 "001000000010110010010101",
						 "001000000010110100110000",
						 "001000000010110111001011",
						 "001000000010111001100110",
						 "001000000010111100000001",
						 "001000000100111010101010",
						 "001000000100111101000101",
						 "001000000100111111100000",
						 "001000000101000001111011",
						 "001000000101000100010110",
						 "001000000101000110110001",
						 "001000000101001001001100",
						 "001000000101001011100111",
						 "001000000101001110000010",
						 "001000000101010000011101",
						 "001000000101010010111000",
						 "001000000101010101010011",
						 "001000000101010111101110",
						 "001000000101011010001001",
						 "001000000101011100100100",
						 "001000000101011110111111",
						 "001000000100111010101010",
						 "001000000100111101000100",
						 "001000000100111111011110",
						 "001000000101000001111000",
						 "001000000101000100010010",
						 "001000000101000110101100",
						 "001000000101001001000110",
						 "001000000101001011100000",
						 "001000000101001101111010",
						 "001000000101010000010100",
						 "001000000101010010101110",
						 "001000000101010101001000",
						 "001000000101010111100010",
						 "001000000101011001111100",
						 "001000000101011100010110",
						 "001000000101011110110000",
						 "001000000100111010101010",
						 "001000000100111101000100",
						 "001000000100111111011110",
						 "001000000101000001111000",
						 "001000000101000100010010",
						 "001000000101000110101100",
						 "001000000101001001000110",
						 "001000000101001011100000",
						 "001000000101001101111010",
						 "001000000101010000010100",
						 "001000000101010010101110",
						 "001000000101010101001000",
						 "001000000101010111100010",
						 "001000000101011001111100",
						 "001000000101011100010110",
						 "001000000101011110110000",
						 "001000000100111010101010",
						 "001000000100111101000100",
						 "001000000100111111011110",
						 "001000000101000001111000",
						 "001000000101000100010010",
						 "001000000101000110101100",
						 "001000000101001001000110",
						 "001000000101001011100000",
						 "001000000101001101111010",
						 "001000000101010000010100",
						 "001000000101010010101110",
						 "001000000101010101001000",
						 "001000000101010111100010",
						 "001000000101011001111100",
						 "001000000101011100010110",
						 "001000000101011110110000",
						 "001000000111011101101000",
						 "001000000111100000000001",
						 "001000000111100010011010",
						 "001000000111100100110011",
						 "001000000111100111001100",
						 "001000000111101001100101",
						 "001000000111101011111110",
						 "001000000111101110010111",
						 "001000000111110000110000",
						 "001000000111110011001001",
						 "001000000111110101100010",
						 "001000000111110111111011",
						 "001000000111111010010100",
						 "001000000111111100101101",
						 "001000000111111111000110",
						 "001000001000000001011111",
						 "001000000111011101101000",
						 "001000000111100000000001",
						 "001000000111100010011010",
						 "001000000111100100110011",
						 "001000000111100111001100",
						 "001000000111101001100101",
						 "001000000111101011111110",
						 "001000000111101110010111",
						 "001000000111110000110000",
						 "001000000111110011001001",
						 "001000000111110101100010",
						 "001000000111110111111011",
						 "001000000111111010010100",
						 "001000000111111100101101",
						 "001000000111111111000110",
						 "001000001000000001011111",
						 "001000000111011101101000",
						 "001000000111100000000001",
						 "001000000111100010011010",
						 "001000000111100100110011",
						 "001000000111100111001100",
						 "001000000111101001100101",
						 "001000000111101011111110",
						 "001000000111101110010111",
						 "001000000111110000110000",
						 "001000000111110011001001",
						 "001000000111110101100010",
						 "001000000111110111111011",
						 "001000000111111010010100",
						 "001000000111111100101101",
						 "001000000111111111000110",
						 "001000001000000001011111",
						 "001000000111011101101000",
						 "001000000111100000000000",
						 "001000000111100010011000",
						 "001000000111100100110000",
						 "001000000111100111001000",
						 "001000000111101001100000",
						 "001000000111101011111000",
						 "001000000111101110010000",
						 "001000000111110000101000",
						 "001000000111110011000000",
						 "001000000111110101011000",
						 "001000000111110111110000",
						 "001000000111111010001000",
						 "001000000111111100100000",
						 "001000000111111110111000",
						 "001000001000000001010000",
						 "001000001010000000100110",
						 "001000001010000010111110",
						 "001000001010000101010110",
						 "001000001010000111101110",
						 "001000001010001010000110",
						 "001000001010001100011110",
						 "001000001010001110110110",
						 "001000001010010001001110",
						 "001000001010010011100110",
						 "001000001010010101111110",
						 "001000001010011000010110",
						 "001000001010011010101110",
						 "001000001010011101000110",
						 "001000001010011111011110",
						 "001000001010100001110110",
						 "001000001010100100001110",
						 "001000001010000000100110",
						 "001000001010000010111110",
						 "001000001010000101010110",
						 "001000001010000111101110",
						 "001000001010001010000110",
						 "001000001010001100011110",
						 "001000001010001110110110",
						 "001000001010010001001110",
						 "001000001010010011100110",
						 "001000001010010101111110",
						 "001000001010011000010110",
						 "001000001010011010101110",
						 "001000001010011101000110",
						 "001000001010011111011110",
						 "001000001010100001110110",
						 "001000001010100100001110",
						 "001000001010000000100110",
						 "001000001010000010111101",
						 "001000001010000101010100",
						 "001000001010000111101011",
						 "001000001010001010000010",
						 "001000001010001100011001",
						 "001000001010001110110000",
						 "001000001010010001000111",
						 "001000001010010011011110",
						 "001000001010010101110101",
						 "001000001010011000001100",
						 "001000001010011010100011",
						 "001000001010011100111010",
						 "001000001010011111010001",
						 "001000001010100001101000",
						 "001000001010100011111111",
						 "001000001010000000100110",
						 "001000001010000010111101",
						 "001000001010000101010100",
						 "001000001010000111101011",
						 "001000001010001010000010",
						 "001000001010001100011001",
						 "001000001010001110110000",
						 "001000001010010001000111",
						 "001000001010010011011110",
						 "001000001010010101110101",
						 "001000001010011000001100",
						 "001000001010011010100011",
						 "001000001010011100111010",
						 "001000001010011111010001",
						 "001000001010100001101000",
						 "001000001010100011111111",
						 "001000001100100011100100",
						 "001000001100100101111011",
						 "001000001100101000010010",
						 "001000001100101010101001",
						 "001000001100101101000000",
						 "001000001100101111010111",
						 "001000001100110001101110",
						 "001000001100110100000101",
						 "001000001100110110011100",
						 "001000001100111000110011",
						 "001000001100111011001010",
						 "001000001100111101100001",
						 "001000001100111111111000",
						 "001000001101000010001111",
						 "001000001101000100100110",
						 "001000001101000110111101",
						 "001000001100100011100100",
						 "001000001100100101111010",
						 "001000001100101000010000",
						 "001000001100101010100110",
						 "001000001100101100111100",
						 "001000001100101111010010",
						 "001000001100110001101000",
						 "001000001100110011111110",
						 "001000001100110110010100",
						 "001000001100111000101010",
						 "001000001100111011000000",
						 "001000001100111101010110",
						 "001000001100111111101100",
						 "001000001101000010000010",
						 "001000001101000100011000",
						 "001000001101000110101110",
						 "001000001100100011100100",
						 "001000001100100101111010",
						 "001000001100101000010000",
						 "001000001100101010100110",
						 "001000001100101100111100",
						 "001000001100101111010010",
						 "001000001100110001101000",
						 "001000001100110011111110",
						 "001000001100110110010100",
						 "001000001100111000101010",
						 "001000001100111011000000",
						 "001000001100111101010110",
						 "001000001100111111101100",
						 "001000001101000010000010",
						 "001000001101000100011000",
						 "001000001101000110101110",
						 "001000001100100011100100",
						 "001000001100100101111010",
						 "001000001100101000010000",
						 "001000001100101010100110",
						 "001000001100101100111100",
						 "001000001100101111010010",
						 "001000001100110001101000",
						 "001000001100110011111110",
						 "001000001100110110010100",
						 "001000001100111000101010",
						 "001000001100111011000000",
						 "001000001100111101010110",
						 "001000001100111111101100",
						 "001000001101000010000010",
						 "001000001101000100011000",
						 "001000001101000110101110",
						 "001000001100100011100100",
						 "001000001100100101111010",
						 "001000001100101000010000",
						 "001000001100101010100110",
						 "001000001100101100111100",
						 "001000001100101111010010",
						 "001000001100110001101000",
						 "001000001100110011111110",
						 "001000001100110110010100",
						 "001000001100111000101010",
						 "001000001100111011000000",
						 "001000001100111101010110",
						 "001000001100111111101100",
						 "001000001101000010000010",
						 "001000001101000100011000",
						 "001000001101000110101110",
						 "001000001111000110100010",
						 "001000001111001000110111",
						 "001000001111001011001100",
						 "001000001111001101100001",
						 "001000001111001111110110",
						 "001000001111010010001011",
						 "001000001111010100100000",
						 "001000001111010110110101",
						 "001000001111011001001010",
						 "001000001111011011011111",
						 "001000001111011101110100",
						 "001000001111100000001001",
						 "001000001111100010011110",
						 "001000001111100100110011",
						 "001000001111100111001000",
						 "001000001111101001011101",
						 "001000001111000110100010",
						 "001000001111001000110111",
						 "001000001111001011001100",
						 "001000001111001101100001",
						 "001000001111001111110110",
						 "001000001111010010001011",
						 "001000001111010100100000",
						 "001000001111010110110101",
						 "001000001111011001001010",
						 "001000001111011011011111",
						 "001000001111011101110100",
						 "001000001111100000001001",
						 "001000001111100010011110",
						 "001000001111100100110011",
						 "001000001111100111001000",
						 "001000001111101001011101",
						 "001000001111000110100010",
						 "001000001111001000110111",
						 "001000001111001011001100",
						 "001000001111001101100001",
						 "001000001111001111110110",
						 "001000001111010010001011",
						 "001000001111010100100000",
						 "001000001111010110110101",
						 "001000001111011001001010",
						 "001000001111011011011111",
						 "001000001111011101110100",
						 "001000001111100000001001",
						 "001000001111100010011110",
						 "001000001111100100110011",
						 "001000001111100111001000",
						 "001000001111101001011101",
						 "001000001111000110100010",
						 "001000001111001000110110",
						 "001000001111001011001010",
						 "001000001111001101011110",
						 "001000001111001111110010",
						 "001000001111010010000110",
						 "001000001111010100011010",
						 "001000001111010110101110",
						 "001000001111011001000010",
						 "001000001111011011010110",
						 "001000001111011101101010",
						 "001000001111011111111110",
						 "001000001111100010010010",
						 "001000001111100100100110",
						 "001000001111100110111010",
						 "001000001111101001001110",
						 "001000010001101001100000",
						 "001000010001101011110100",
						 "001000010001101110001000",
						 "001000010001110000011100",
						 "001000010001110010110000",
						 "001000010001110101000100",
						 "001000010001110111011000",
						 "001000010001111001101100",
						 "001000010001111100000000",
						 "001000010001111110010100",
						 "001000010010000000101000",
						 "001000010010000010111100",
						 "001000010010000101010000",
						 "001000010010000111100100",
						 "001000010010001001111000",
						 "001000010010001100001100",
						 "001000010001101001100000",
						 "001000010001101011110100",
						 "001000010001101110001000",
						 "001000010001110000011100",
						 "001000010001110010110000",
						 "001000010001110101000100",
						 "001000010001110111011000",
						 "001000010001111001101100",
						 "001000010001111100000000",
						 "001000010001111110010100",
						 "001000010010000000101000",
						 "001000010010000010111100",
						 "001000010010000101010000",
						 "001000010010000111100100",
						 "001000010010001001111000",
						 "001000010010001100001100",
						 "001000010001101001100000",
						 "001000010001101011110011",
						 "001000010001101110000110",
						 "001000010001110000011001",
						 "001000010001110010101100",
						 "001000010001110100111111",
						 "001000010001110111010010",
						 "001000010001111001100101",
						 "001000010001111011111000",
						 "001000010001111110001011",
						 "001000010010000000011110",
						 "001000010010000010110001",
						 "001000010010000101000100",
						 "001000010010000111010111",
						 "001000010010001001101010",
						 "001000010010001011111101",
						 "001000010001101001100000",
						 "001000010001101011110011",
						 "001000010001101110000110",
						 "001000010001110000011001",
						 "001000010001110010101100",
						 "001000010001110100111111",
						 "001000010001110111010010",
						 "001000010001111001100101",
						 "001000010001111011111000",
						 "001000010001111110001011",
						 "001000010010000000011110",
						 "001000010010000010110001",
						 "001000010010000101000100",
						 "001000010010000111010111",
						 "001000010010001001101010",
						 "001000010010001011111101",
						 "001000010001101001100000",
						 "001000010001101011110011",
						 "001000010001101110000110",
						 "001000010001110000011001",
						 "001000010001110010101100",
						 "001000010001110100111111",
						 "001000010001110111010010",
						 "001000010001111001100101",
						 "001000010001111011111000",
						 "001000010001111110001011",
						 "001000010010000000011110",
						 "001000010010000010110001",
						 "001000010010000101000100",
						 "001000010010000111010111",
						 "001000010010001001101010",
						 "001000010010001011111101",
						 "001000010100001100011110",
						 "001000010100001110110000",
						 "001000010100010001000010",
						 "001000010100010011010100",
						 "001000010100010101100110",
						 "001000010100010111111000",
						 "001000010100011010001010",
						 "001000010100011100011100",
						 "001000010100011110101110",
						 "001000010100100001000000",
						 "001000010100100011010010",
						 "001000010100100101100100",
						 "001000010100100111110110",
						 "001000010100101010001000",
						 "001000010100101100011010",
						 "001000010100101110101100",
						 "001000010100001100011110",
						 "001000010100001110110000",
						 "001000010100010001000010",
						 "001000010100010011010100",
						 "001000010100010101100110",
						 "001000010100010111111000",
						 "001000010100011010001010",
						 "001000010100011100011100",
						 "001000010100011110101110",
						 "001000010100100001000000",
						 "001000010100100011010010",
						 "001000010100100101100100",
						 "001000010100100111110110",
						 "001000010100101010001000",
						 "001000010100101100011010",
						 "001000010100101110101100",
						 "001000010100001100011110",
						 "001000010100001110110000",
						 "001000010100010001000010",
						 "001000010100010011010100",
						 "001000010100010101100110",
						 "001000010100010111111000",
						 "001000010100011010001010",
						 "001000010100011100011100",
						 "001000010100011110101110",
						 "001000010100100001000000",
						 "001000010100100011010010",
						 "001000010100100101100100",
						 "001000010100100111110110",
						 "001000010100101010001000",
						 "001000010100101100011010",
						 "001000010100101110101100",
						 "001000010100001100011110",
						 "001000010100001110101111",
						 "001000010100010001000000",
						 "001000010100010011010001",
						 "001000010100010101100010",
						 "001000010100010111110011",
						 "001000010100011010000100",
						 "001000010100011100010101",
						 "001000010100011110100110",
						 "001000010100100000110111",
						 "001000010100100011001000",
						 "001000010100100101011001",
						 "001000010100100111101010",
						 "001000010100101001111011",
						 "001000010100101100001100",
						 "001000010100101110011101",
						 "001000010110101111011100",
						 "001000010110110001101101",
						 "001000010110110011111110",
						 "001000010110110110001111",
						 "001000010110111000100000",
						 "001000010110111010110001",
						 "001000010110111101000010",
						 "001000010110111111010011",
						 "001000010111000001100100",
						 "001000010111000011110101",
						 "001000010111000110000110",
						 "001000010111001000010111",
						 "001000010111001010101000",
						 "001000010111001100111001",
						 "001000010111001111001010",
						 "001000010111010001011011",
						 "001000010110101111011100",
						 "001000010110110001101101",
						 "001000010110110011111110",
						 "001000010110110110001111",
						 "001000010110111000100000",
						 "001000010110111010110001",
						 "001000010110111101000010",
						 "001000010110111111010011",
						 "001000010111000001100100",
						 "001000010111000011110101",
						 "001000010111000110000110",
						 "001000010111001000010111",
						 "001000010111001010101000",
						 "001000010111001100111001",
						 "001000010111001111001010",
						 "001000010111010001011011",
						 "001000010110101111011100",
						 "001000010110110001101100",
						 "001000010110110011111100",
						 "001000010110110110001100",
						 "001000010110111000011100",
						 "001000010110111010101100",
						 "001000010110111100111100",
						 "001000010110111111001100",
						 "001000010111000001011100",
						 "001000010111000011101100",
						 "001000010111000101111100",
						 "001000010111001000001100",
						 "001000010111001010011100",
						 "001000010111001100101100",
						 "001000010111001110111100",
						 "001000010111010001001100",
						 "001000010110101111011100",
						 "001000010110110001101100",
						 "001000010110110011111100",
						 "001000010110110110001100",
						 "001000010110111000011100",
						 "001000010110111010101100",
						 "001000010110111100111100",
						 "001000010110111111001100",
						 "001000010111000001011100",
						 "001000010111000011101100",
						 "001000010111000101111100",
						 "001000010111001000001100",
						 "001000010111001010011100",
						 "001000010111001100101100",
						 "001000010111001110111100",
						 "001000010111010001001100",
						 "001000010110101111011100",
						 "001000010110110001101100",
						 "001000010110110011111100",
						 "001000010110110110001100",
						 "001000010110111000011100",
						 "001000010110111010101100",
						 "001000010110111100111100",
						 "001000010110111111001100",
						 "001000010111000001011100",
						 "001000010111000011101100",
						 "001000010111000101111100",
						 "001000010111001000001100",
						 "001000010111001010011100",
						 "001000010111001100101100",
						 "001000010111001110111100",
						 "001000010111010001001100",
						 "001000011001010010011010",
						 "001000011001010100101001",
						 "001000011001010110111000",
						 "001000011001011001000111",
						 "001000011001011011010110",
						 "001000011001011101100101",
						 "001000011001011111110100",
						 "001000011001100010000011",
						 "001000011001100100010010",
						 "001000011001100110100001",
						 "001000011001101000110000",
						 "001000011001101010111111",
						 "001000011001101101001110",
						 "001000011001101111011101",
						 "001000011001110001101100",
						 "001000011001110011111011",
						 "001000011001010010011010",
						 "001000011001010100101001",
						 "001000011001010110111000",
						 "001000011001011001000111",
						 "001000011001011011010110",
						 "001000011001011101100101",
						 "001000011001011111110100",
						 "001000011001100010000011",
						 "001000011001100100010010",
						 "001000011001100110100001",
						 "001000011001101000110000",
						 "001000011001101010111111",
						 "001000011001101101001110",
						 "001000011001101111011101",
						 "001000011001110001101100",
						 "001000011001110011111011",
						 "001000011001010010011010",
						 "001000011001010100101001",
						 "001000011001010110111000",
						 "001000011001011001000111",
						 "001000011001011011010110",
						 "001000011001011101100101",
						 "001000011001011111110100",
						 "001000011001100010000011",
						 "001000011001100100010010",
						 "001000011001100110100001",
						 "001000011001101000110000",
						 "001000011001101010111111",
						 "001000011001101101001110",
						 "001000011001101111011101",
						 "001000011001110001101100",
						 "001000011001110011111011",
						 "001000011001010010011010",
						 "001000011001010100101000",
						 "001000011001010110110110",
						 "001000011001011001000100",
						 "001000011001011011010010",
						 "001000011001011101100000",
						 "001000011001011111101110",
						 "001000011001100001111100",
						 "001000011001100100001010",
						 "001000011001100110011000",
						 "001000011001101000100110",
						 "001000011001101010110100",
						 "001000011001101101000010",
						 "001000011001101111010000",
						 "001000011001110001011110",
						 "001000011001110011101100",
						 "001000011011110101011000",
						 "001000011011110111100110",
						 "001000011011111001110100",
						 "001000011011111100000010",
						 "001000011011111110010000",
						 "001000011100000000011110",
						 "001000011100000010101100",
						 "001000011100000100111010",
						 "001000011100000111001000",
						 "001000011100001001010110",
						 "001000011100001011100100",
						 "001000011100001101110010",
						 "001000011100010000000000",
						 "001000011100010010001110",
						 "001000011100010100011100",
						 "001000011100010110101010",
						 "001000011011110101011000",
						 "001000011011110111100110",
						 "001000011011111001110100",
						 "001000011011111100000010",
						 "001000011011111110010000",
						 "001000011100000000011110",
						 "001000011100000010101100",
						 "001000011100000100111010",
						 "001000011100000111001000",
						 "001000011100001001010110",
						 "001000011100001011100100",
						 "001000011100001101110010",
						 "001000011100010000000000",
						 "001000011100010010001110",
						 "001000011100010100011100",
						 "001000011100010110101010",
						 "001000011011110101011000",
						 "001000011011110111100110",
						 "001000011011111001110100",
						 "001000011011111100000010",
						 "001000011011111110010000",
						 "001000011100000000011110",
						 "001000011100000010101100",
						 "001000011100000100111010",
						 "001000011100000111001000",
						 "001000011100001001010110",
						 "001000011100001011100100",
						 "001000011100001101110010",
						 "001000011100010000000000",
						 "001000011100010010001110",
						 "001000011100010100011100",
						 "001000011100010110101010",
						 "001000011011110101011000",
						 "001000011011110111100101",
						 "001000011011111001110010",
						 "001000011011111011111111",
						 "001000011011111110001100",
						 "001000011100000000011001",
						 "001000011100000010100110",
						 "001000011100000100110011",
						 "001000011100000111000000",
						 "001000011100001001001101",
						 "001000011100001011011010",
						 "001000011100001101100111",
						 "001000011100001111110100",
						 "001000011100010010000001",
						 "001000011100010100001110",
						 "001000011100010110011011",
						 "001000011011110101011000",
						 "001000011011110111100101",
						 "001000011011111001110010",
						 "001000011011111011111111",
						 "001000011011111110001100",
						 "001000011100000000011001",
						 "001000011100000010100110",
						 "001000011100000100110011",
						 "001000011100000111000000",
						 "001000011100001001001101",
						 "001000011100001011011010",
						 "001000011100001101100111",
						 "001000011100001111110100",
						 "001000011100010010000001",
						 "001000011100010100001110",
						 "001000011100010110011011",
						 "001000011110011000010110",
						 "001000011110011010100011",
						 "001000011110011100110000",
						 "001000011110011110111101",
						 "001000011110100001001010",
						 "001000011110100011010111",
						 "001000011110100101100100",
						 "001000011110100111110001",
						 "001000011110101001111110",
						 "001000011110101100001011",
						 "001000011110101110011000",
						 "001000011110110000100101",
						 "001000011110110010110010",
						 "001000011110110100111111",
						 "001000011110110111001100",
						 "001000011110111001011001",
						 "001000011110011000010110",
						 "001000011110011010100010",
						 "001000011110011100101110",
						 "001000011110011110111010",
						 "001000011110100001000110",
						 "001000011110100011010010",
						 "001000011110100101011110",
						 "001000011110100111101010",
						 "001000011110101001110110",
						 "001000011110101100000010",
						 "001000011110101110001110",
						 "001000011110110000011010",
						 "001000011110110010100110",
						 "001000011110110100110010",
						 "001000011110110110111110",
						 "001000011110111001001010",
						 "001000011110011000010110",
						 "001000011110011010100010",
						 "001000011110011100101110",
						 "001000011110011110111010",
						 "001000011110100001000110",
						 "001000011110100011010010",
						 "001000011110100101011110",
						 "001000011110100111101010",
						 "001000011110101001110110",
						 "001000011110101100000010",
						 "001000011110101110001110",
						 "001000011110110000011010",
						 "001000011110110010100110",
						 "001000011110110100110010",
						 "001000011110110110111110",
						 "001000011110111001001010",
						 "001000011110011000010110",
						 "001000011110011010100010",
						 "001000011110011100101110",
						 "001000011110011110111010",
						 "001000011110100001000110",
						 "001000011110100011010010",
						 "001000011110100101011110",
						 "001000011110100111101010",
						 "001000011110101001110110",
						 "001000011110101100000010",
						 "001000011110101110001110",
						 "001000011110110000011010",
						 "001000011110110010100110",
						 "001000011110110100110010",
						 "001000011110110110111110",
						 "001000011110111001001010",
						 "001000100000111011010100",
						 "001000100000111101011111",
						 "001000100000111111101010",
						 "001000100001000001110101",
						 "001000100001000100000000",
						 "001000100001000110001011",
						 "001000100001001000010110",
						 "001000100001001010100001",
						 "001000100001001100101100",
						 "001000100001001110110111",
						 "001000100001010001000010",
						 "001000100001010011001101",
						 "001000100001010101011000",
						 "001000100001010111100011",
						 "001000100001011001101110",
						 "001000100001011011111001",
						 "001000100000111011010100",
						 "001000100000111101011111",
						 "001000100000111111101010",
						 "001000100001000001110101",
						 "001000100001000100000000",
						 "001000100001000110001011",
						 "001000100001001000010110",
						 "001000100001001010100001",
						 "001000100001001100101100",
						 "001000100001001110110111",
						 "001000100001010001000010",
						 "001000100001010011001101",
						 "001000100001010101011000",
						 "001000100001010111100011",
						 "001000100001011001101110",
						 "001000100001011011111001",
						 "001000100000111011010100",
						 "001000100000111101011111",
						 "001000100000111111101010",
						 "001000100001000001110101",
						 "001000100001000100000000",
						 "001000100001000110001011",
						 "001000100001001000010110",
						 "001000100001001010100001",
						 "001000100001001100101100",
						 "001000100001001110110111",
						 "001000100001010001000010",
						 "001000100001010011001101",
						 "001000100001010101011000",
						 "001000100001010111100011",
						 "001000100001011001101110",
						 "001000100001011011111001",
						 "001000100000111011010100",
						 "001000100000111101011110",
						 "001000100000111111101000",
						 "001000100001000001110010",
						 "001000100001000011111100",
						 "001000100001000110000110",
						 "001000100001001000010000",
						 "001000100001001010011010",
						 "001000100001001100100100",
						 "001000100001001110101110",
						 "001000100001010000111000",
						 "001000100001010011000010",
						 "001000100001010101001100",
						 "001000100001010111010110",
						 "001000100001011001100000",
						 "001000100001011011101010",
						 "001000100000111011010100",
						 "001000100000111101011110",
						 "001000100000111111101000",
						 "001000100001000001110010",
						 "001000100001000011111100",
						 "001000100001000110000110",
						 "001000100001001000010000",
						 "001000100001001010011010",
						 "001000100001001100100100",
						 "001000100001001110101110",
						 "001000100001010000111000",
						 "001000100001010011000010",
						 "001000100001010101001100",
						 "001000100001010111010110",
						 "001000100001011001100000",
						 "001000100001011011101010",
						 "001000100011011110010010",
						 "001000100011100000011100",
						 "001000100011100010100110",
						 "001000100011100100110000",
						 "001000100011100110111010",
						 "001000100011101001000100",
						 "001000100011101011001110",
						 "001000100011101101011000",
						 "001000100011101111100010",
						 "001000100011110001101100",
						 "001000100011110011110110",
						 "001000100011110110000000",
						 "001000100011111000001010",
						 "001000100011111010010100",
						 "001000100011111100011110",
						 "001000100011111110101000",
						 "001000100011011110010010",
						 "001000100011100000011011",
						 "001000100011100010100100",
						 "001000100011100100101101",
						 "001000100011100110110110",
						 "001000100011101000111111",
						 "001000100011101011001000",
						 "001000100011101101010001",
						 "001000100011101111011010",
						 "001000100011110001100011",
						 "001000100011110011101100",
						 "001000100011110101110101",
						 "001000100011110111111110",
						 "001000100011111010000111",
						 "001000100011111100010000",
						 "001000100011111110011001",
						 "001000100011011110010010",
						 "001000100011100000011011",
						 "001000100011100010100100",
						 "001000100011100100101101",
						 "001000100011100110110110",
						 "001000100011101000111111",
						 "001000100011101011001000",
						 "001000100011101101010001",
						 "001000100011101111011010",
						 "001000100011110001100011",
						 "001000100011110011101100",
						 "001000100011110101110101",
						 "001000100011110111111110",
						 "001000100011111010000111",
						 "001000100011111100010000",
						 "001000100011111110011001",
						 "001000100011011110010010",
						 "001000100011100000011011",
						 "001000100011100010100100",
						 "001000100011100100101101",
						 "001000100011100110110110",
						 "001000100011101000111111",
						 "001000100011101011001000",
						 "001000100011101101010001",
						 "001000100011101111011010",
						 "001000100011110001100011",
						 "001000100011110011101100",
						 "001000100011110101110101",
						 "001000100011110111111110",
						 "001000100011111010000111",
						 "001000100011111100010000",
						 "001000100011111110011001",
						 "001000100011011110010010",
						 "001000100011100000011010",
						 "001000100011100010100010",
						 "001000100011100100101010",
						 "001000100011100110110010",
						 "001000100011101000111010",
						 "001000100011101011000010",
						 "001000100011101101001010",
						 "001000100011101111010010",
						 "001000100011110001011010",
						 "001000100011110011100010",
						 "001000100011110101101010",
						 "001000100011110111110010",
						 "001000100011111001111010",
						 "001000100011111100000010",
						 "001000100011111110001010",
						 "001000100110000001010000",
						 "001000100110000011011000",
						 "001000100110000101100000",
						 "001000100110000111101000",
						 "001000100110001001110000",
						 "001000100110001011111000",
						 "001000100110001110000000",
						 "001000100110010000001000",
						 "001000100110010010010000",
						 "001000100110010100011000",
						 "001000100110010110100000",
						 "001000100110011000101000",
						 "001000100110011010110000",
						 "001000100110011100111000",
						 "001000100110011111000000",
						 "001000100110100001001000",
						 "001000100110000001010000",
						 "001000100110000011011000",
						 "001000100110000101100000",
						 "001000100110000111101000",
						 "001000100110001001110000",
						 "001000100110001011111000",
						 "001000100110001110000000",
						 "001000100110010000001000",
						 "001000100110010010010000",
						 "001000100110010100011000",
						 "001000100110010110100000",
						 "001000100110011000101000",
						 "001000100110011010110000",
						 "001000100110011100111000",
						 "001000100110011111000000",
						 "001000100110100001001000",
						 "001000100110000001010000",
						 "001000100110000011010111",
						 "001000100110000101011110",
						 "001000100110000111100101",
						 "001000100110001001101100",
						 "001000100110001011110011",
						 "001000100110001101111010",
						 "001000100110010000000001",
						 "001000100110010010001000",
						 "001000100110010100001111",
						 "001000100110010110010110",
						 "001000100110011000011101",
						 "001000100110011010100100",
						 "001000100110011100101011",
						 "001000100110011110110010",
						 "001000100110100000111001",
						 "001000100110000001010000",
						 "001000100110000011010111",
						 "001000100110000101011110",
						 "001000100110000111100101",
						 "001000100110001001101100",
						 "001000100110001011110011",
						 "001000100110001101111010",
						 "001000100110010000000001",
						 "001000100110010010001000",
						 "001000100110010100001111",
						 "001000100110010110010110",
						 "001000100110011000011101",
						 "001000100110011010100100",
						 "001000100110011100101011",
						 "001000100110011110110010",
						 "001000100110100000111001",
						 "001000100110000001010000",
						 "001000100110000011010111",
						 "001000100110000101011110",
						 "001000100110000111100101",
						 "001000100110001001101100",
						 "001000100110001011110011",
						 "001000100110001101111010",
						 "001000100110010000000001",
						 "001000100110010010001000",
						 "001000100110010100001111",
						 "001000100110010110010110",
						 "001000100110011000011101",
						 "001000100110011010100100",
						 "001000100110011100101011",
						 "001000100110011110110010",
						 "001000100110100000111001",
						 "001000101000100100001110",
						 "001000101000100110010100",
						 "001000101000101000011010",
						 "001000101000101010100000",
						 "001000101000101100100110",
						 "001000101000101110101100",
						 "001000101000110000110010",
						 "001000101000110010111000",
						 "001000101000110100111110",
						 "001000101000110111000100",
						 "001000101000111001001010",
						 "001000101000111011010000",
						 "001000101000111101010110",
						 "001000101000111111011100",
						 "001000101001000001100010",
						 "001000101001000011101000",
						 "001000101000100100001110",
						 "001000101000100110010100",
						 "001000101000101000011010",
						 "001000101000101010100000",
						 "001000101000101100100110",
						 "001000101000101110101100",
						 "001000101000110000110010",
						 "001000101000110010111000",
						 "001000101000110100111110",
						 "001000101000110111000100",
						 "001000101000111001001010",
						 "001000101000111011010000",
						 "001000101000111101010110",
						 "001000101000111111011100",
						 "001000101001000001100010",
						 "001000101001000011101000",
						 "001000101000100100001110",
						 "001000101000100110010100",
						 "001000101000101000011010",
						 "001000101000101010100000",
						 "001000101000101100100110",
						 "001000101000101110101100",
						 "001000101000110000110010",
						 "001000101000110010111000",
						 "001000101000110100111110",
						 "001000101000110111000100",
						 "001000101000111001001010",
						 "001000101000111011010000",
						 "001000101000111101010110",
						 "001000101000111111011100",
						 "001000101001000001100010",
						 "001000101001000011101000",
						 "001000101000100100001110",
						 "001000101000100110010011",
						 "001000101000101000011000",
						 "001000101000101010011101",
						 "001000101000101100100010",
						 "001000101000101110100111",
						 "001000101000110000101100",
						 "001000101000110010110001",
						 "001000101000110100110110",
						 "001000101000110110111011",
						 "001000101000111001000000",
						 "001000101000111011000101",
						 "001000101000111101001010",
						 "001000101000111111001111",
						 "001000101001000001010100",
						 "001000101001000011011001",
						 "001000101011000111001100",
						 "001000101011001001010001",
						 "001000101011001011010110",
						 "001000101011001101011011",
						 "001000101011001111100000",
						 "001000101011010001100101",
						 "001000101011010011101010",
						 "001000101011010101101111",
						 "001000101011010111110100",
						 "001000101011011001111001",
						 "001000101011011011111110",
						 "001000101011011110000011",
						 "001000101011100000001000",
						 "001000101011100010001101",
						 "001000101011100100010010",
						 "001000101011100110010111",
						 "001000101011000111001100",
						 "001000101011001001010001",
						 "001000101011001011010110",
						 "001000101011001101011011",
						 "001000101011001111100000",
						 "001000101011010001100101",
						 "001000101011010011101010",
						 "001000101011010101101111",
						 "001000101011010111110100",
						 "001000101011011001111001",
						 "001000101011011011111110",
						 "001000101011011110000011",
						 "001000101011100000001000",
						 "001000101011100010001101",
						 "001000101011100100010010",
						 "001000101011100110010111",
						 "001000101011000111001100",
						 "001000101011001001010000",
						 "001000101011001011010100",
						 "001000101011001101011000",
						 "001000101011001111011100",
						 "001000101011010001100000",
						 "001000101011010011100100",
						 "001000101011010101101000",
						 "001000101011010111101100",
						 "001000101011011001110000",
						 "001000101011011011110100",
						 "001000101011011101111000",
						 "001000101011011111111100",
						 "001000101011100010000000",
						 "001000101011100100000100",
						 "001000101011100110001000",
						 "001000101011000111001100",
						 "001000101011001001010000",
						 "001000101011001011010100",
						 "001000101011001101011000",
						 "001000101011001111011100",
						 "001000101011010001100000",
						 "001000101011010011100100",
						 "001000101011010101101000",
						 "001000101011010111101100",
						 "001000101011011001110000",
						 "001000101011011011110100",
						 "001000101011011101111000",
						 "001000101011011111111100",
						 "001000101011100010000000",
						 "001000101011100100000100",
						 "001000101011100110001000",
						 "001000101011000111001100",
						 "001000101011001001010000",
						 "001000101011001011010100",
						 "001000101011001101011000",
						 "001000101011001111011100",
						 "001000101011010001100000",
						 "001000101011010011100100",
						 "001000101011010101101000",
						 "001000101011010111101100",
						 "001000101011011001110000",
						 "001000101011011011110100",
						 "001000101011011101111000",
						 "001000101011011111111100",
						 "001000101011100010000000",
						 "001000101011100100000100",
						 "001000101011100110001000",
						 "001000101101101010001010",
						 "001000101101101100001101",
						 "001000101101101110010000",
						 "001000101101110000010011",
						 "001000101101110010010110",
						 "001000101101110100011001",
						 "001000101101110110011100",
						 "001000101101111000011111",
						 "001000101101111010100010",
						 "001000101101111100100101",
						 "001000101101111110101000",
						 "001000101110000000101011",
						 "001000101110000010101110",
						 "001000101110000100110001",
						 "001000101110000110110100",
						 "001000101110001000110111",
						 "001000101101101010001010",
						 "001000101101101100001101",
						 "001000101101101110010000",
						 "001000101101110000010011",
						 "001000101101110010010110",
						 "001000101101110100011001",
						 "001000101101110110011100",
						 "001000101101111000011111",
						 "001000101101111010100010",
						 "001000101101111100100101",
						 "001000101101111110101000",
						 "001000101110000000101011",
						 "001000101110000010101110",
						 "001000101110000100110001",
						 "001000101110000110110100",
						 "001000101110001000110111",
						 "001000101101101010001010",
						 "001000101101101100001101",
						 "001000101101101110010000",
						 "001000101101110000010011",
						 "001000101101110010010110",
						 "001000101101110100011001",
						 "001000101101110110011100",
						 "001000101101111000011111",
						 "001000101101111010100010",
						 "001000101101111100100101",
						 "001000101101111110101000",
						 "001000101110000000101011",
						 "001000101110000010101110",
						 "001000101110000100110001",
						 "001000101110000110110100",
						 "001000101110001000110111",
						 "001000101101101010001010",
						 "001000101101101100001100",
						 "001000101101101110001110",
						 "001000101101110000010000",
						 "001000101101110010010010",
						 "001000101101110100010100",
						 "001000101101110110010110",
						 "001000101101111000011000",
						 "001000101101111010011010",
						 "001000101101111100011100",
						 "001000101101111110011110",
						 "001000101110000000100000",
						 "001000101110000010100010",
						 "001000101110000100100100",
						 "001000101110000110100110",
						 "001000101110001000101000",
						 "001000101101101010001010",
						 "001000101101101100001100",
						 "001000101101101110001110",
						 "001000101101110000010000",
						 "001000101101110010010010",
						 "001000101101110100010100",
						 "001000101101110110010110",
						 "001000101101111000011000",
						 "001000101101111010011010",
						 "001000101101111100011100",
						 "001000101101111110011110",
						 "001000101110000000100000",
						 "001000101110000010100010",
						 "001000101110000100100100",
						 "001000101110000110100110",
						 "001000101110001000101000",
						 "001000110000001101001000",
						 "001000110000001111001010",
						 "001000110000010001001100",
						 "001000110000010011001110",
						 "001000110000010101010000",
						 "001000110000010111010010",
						 "001000110000011001010100",
						 "001000110000011011010110",
						 "001000110000011101011000",
						 "001000110000011111011010",
						 "001000110000100001011100",
						 "001000110000100011011110",
						 "001000110000100101100000",
						 "001000110000100111100010",
						 "001000110000101001100100",
						 "001000110000101011100110",
						 "001000110000001101001000",
						 "001000110000001111001001",
						 "001000110000010001001010",
						 "001000110000010011001011",
						 "001000110000010101001100",
						 "001000110000010111001101",
						 "001000110000011001001110",
						 "001000110000011011001111",
						 "001000110000011101010000",
						 "001000110000011111010001",
						 "001000110000100001010010",
						 "001000110000100011010011",
						 "001000110000100101010100",
						 "001000110000100111010101",
						 "001000110000101001010110",
						 "001000110000101011010111",
						 "001000110000001101001000",
						 "001000110000001111001001",
						 "001000110000010001001010",
						 "001000110000010011001011",
						 "001000110000010101001100",
						 "001000110000010111001101",
						 "001000110000011001001110",
						 "001000110000011011001111",
						 "001000110000011101010000",
						 "001000110000011111010001",
						 "001000110000100001010010",
						 "001000110000100011010011",
						 "001000110000100101010100",
						 "001000110000100111010101",
						 "001000110000101001010110",
						 "001000110000101011010111",
						 "001000110000001101001000",
						 "001000110000001111001001",
						 "001000110000010001001010",
						 "001000110000010011001011",
						 "001000110000010101001100",
						 "001000110000010111001101",
						 "001000110000011001001110",
						 "001000110000011011001111",
						 "001000110000011101010000",
						 "001000110000011111010001",
						 "001000110000100001010010",
						 "001000110000100011010011",
						 "001000110000100101010100",
						 "001000110000100111010101",
						 "001000110000101001010110",
						 "001000110000101011010111",
						 "001000110000001101001000",
						 "001000110000001111001000",
						 "001000110000010001001000",
						 "001000110000010011001000",
						 "001000110000010101001000",
						 "001000110000010111001000",
						 "001000110000011001001000",
						 "001000110000011011001000",
						 "001000110000011101001000",
						 "001000110000011111001000",
						 "001000110000100001001000",
						 "001000110000100011001000",
						 "001000110000100101001000",
						 "001000110000100111001000",
						 "001000110000101001001000",
						 "001000110000101011001000",
						 "001000110010110000000110",
						 "001000110010110010000110",
						 "001000110010110100000110",
						 "001000110010110110000110",
						 "001000110010111000000110",
						 "001000110010111010000110",
						 "001000110010111100000110",
						 "001000110010111110000110",
						 "001000110011000000000110",
						 "001000110011000010000110",
						 "001000110011000100000110",
						 "001000110011000110000110",
						 "001000110011001000000110",
						 "001000110011001010000110",
						 "001000110011001100000110",
						 "001000110011001110000110",
						 "001000110010110000000110",
						 "001000110010110010000110",
						 "001000110010110100000110",
						 "001000110010110110000110",
						 "001000110010111000000110",
						 "001000110010111010000110",
						 "001000110010111100000110",
						 "001000110010111110000110",
						 "001000110011000000000110",
						 "001000110011000010000110",
						 "001000110011000100000110",
						 "001000110011000110000110",
						 "001000110011001000000110",
						 "001000110011001010000110",
						 "001000110011001100000110",
						 "001000110011001110000110",
						 "001000110010110000000110",
						 "001000110010110010000101",
						 "001000110010110100000100",
						 "001000110010110110000011",
						 "001000110010111000000010",
						 "001000110010111010000001",
						 "001000110010111100000000",
						 "001000110010111101111111",
						 "001000110010111111111110",
						 "001000110011000001111101",
						 "001000110011000011111100",
						 "001000110011000101111011",
						 "001000110011000111111010",
						 "001000110011001001111001",
						 "001000110011001011111000",
						 "001000110011001101110111",
						 "001000110010110000000110",
						 "001000110010110010000101",
						 "001000110010110100000100",
						 "001000110010110110000011",
						 "001000110010111000000010",
						 "001000110010111010000001",
						 "001000110010111100000000",
						 "001000110010111101111111",
						 "001000110010111111111110",
						 "001000110011000001111101",
						 "001000110011000011111100",
						 "001000110011000101111011",
						 "001000110011000111111010",
						 "001000110011001001111001",
						 "001000110011001011111000",
						 "001000110011001101110111",
						 "001000110010110000000110",
						 "001000110010110010000101",
						 "001000110010110100000100",
						 "001000110010110110000011",
						 "001000110010111000000010",
						 "001000110010111010000001",
						 "001000110010111100000000",
						 "001000110010111101111111",
						 "001000110010111111111110",
						 "001000110011000001111101",
						 "001000110011000011111100",
						 "001000110011000101111011",
						 "001000110011000111111010",
						 "001000110011001001111001",
						 "001000110011001011111000",
						 "001000110011001101110111",
						 "001000110010110000000110",
						 "001000110010110010000100",
						 "001000110010110100000010",
						 "001000110010110110000000",
						 "001000110010110111111110",
						 "001000110010111001111100",
						 "001000110010111011111010",
						 "001000110010111101111000",
						 "001000110010111111110110",
						 "001000110011000001110100",
						 "001000110011000011110010",
						 "001000110011000101110000",
						 "001000110011000111101110",
						 "001000110011001001101100",
						 "001000110011001011101010",
						 "001000110011001101101000",
						 "001000110101010011000100",
						 "001000110101010101000010",
						 "001000110101010111000000",
						 "001000110101011000111110",
						 "001000110101011010111100",
						 "001000110101011100111010",
						 "001000110101011110111000",
						 "001000110101100000110110",
						 "001000110101100010110100",
						 "001000110101100100110010",
						 "001000110101100110110000",
						 "001000110101101000101110",
						 "001000110101101010101100",
						 "001000110101101100101010",
						 "001000110101101110101000",
						 "001000110101110000100110",
						 "001000110101010011000100",
						 "001000110101010101000010",
						 "001000110101010111000000",
						 "001000110101011000111110",
						 "001000110101011010111100",
						 "001000110101011100111010",
						 "001000110101011110111000",
						 "001000110101100000110110",
						 "001000110101100010110100",
						 "001000110101100100110010",
						 "001000110101100110110000",
						 "001000110101101000101110",
						 "001000110101101010101100",
						 "001000110101101100101010",
						 "001000110101101110101000",
						 "001000110101110000100110",
						 "001000110101010011000100",
						 "001000110101010101000001",
						 "001000110101010110111110",
						 "001000110101011000111011",
						 "001000110101011010111000",
						 "001000110101011100110101",
						 "001000110101011110110010",
						 "001000110101100000101111",
						 "001000110101100010101100",
						 "001000110101100100101001",
						 "001000110101100110100110",
						 "001000110101101000100011",
						 "001000110101101010100000",
						 "001000110101101100011101",
						 "001000110101101110011010",
						 "001000110101110000010111",
						 "001000110101010011000100",
						 "001000110101010101000001",
						 "001000110101010110111110",
						 "001000110101011000111011",
						 "001000110101011010111000",
						 "001000110101011100110101",
						 "001000110101011110110010",
						 "001000110101100000101111",
						 "001000110101100010101100",
						 "001000110101100100101001",
						 "001000110101100110100110",
						 "001000110101101000100011",
						 "001000110101101010100000",
						 "001000110101101100011101",
						 "001000110101101110011010",
						 "001000110101110000010111",
						 "001000110101010011000100",
						 "001000110101010101000000",
						 "001000110101010110111100",
						 "001000110101011000111000",
						 "001000110101011010110100",
						 "001000110101011100110000",
						 "001000110101011110101100",
						 "001000110101100000101000",
						 "001000110101100010100100",
						 "001000110101100100100000",
						 "001000110101100110011100",
						 "001000110101101000011000",
						 "001000110101101010010100",
						 "001000110101101100010000",
						 "001000110101101110001100",
						 "001000110101110000001000",
						 "001000110111110110000010",
						 "001000110111110111111110",
						 "001000110111111001111010",
						 "001000110111111011110110",
						 "001000110111111101110010",
						 "001000110111111111101110",
						 "001000111000000001101010",
						 "001000111000000011100110",
						 "001000111000000101100010",
						 "001000111000000111011110",
						 "001000111000001001011010",
						 "001000111000001011010110",
						 "001000111000001101010010",
						 "001000111000001111001110",
						 "001000111000010001001010",
						 "001000111000010011000110",
						 "001000110111110110000010",
						 "001000110111110111111110",
						 "001000110111111001111010",
						 "001000110111111011110110",
						 "001000110111111101110010",
						 "001000110111111111101110",
						 "001000111000000001101010",
						 "001000111000000011100110",
						 "001000111000000101100010",
						 "001000111000000111011110",
						 "001000111000001001011010",
						 "001000111000001011010110",
						 "001000111000001101010010",
						 "001000111000001111001110",
						 "001000111000010001001010",
						 "001000111000010011000110",
						 "001000110111110110000010",
						 "001000110111110111111101",
						 "001000110111111001111000",
						 "001000110111111011110011",
						 "001000110111111101101110",
						 "001000110111111111101001",
						 "001000111000000001100100",
						 "001000111000000011011111",
						 "001000111000000101011010",
						 "001000111000000111010101",
						 "001000111000001001010000",
						 "001000111000001011001011",
						 "001000111000001101000110",
						 "001000111000001111000001",
						 "001000111000010000111100",
						 "001000111000010010110111",
						 "001000110111110110000010",
						 "001000110111110111111101",
						 "001000110111111001111000",
						 "001000110111111011110011",
						 "001000110111111101101110",
						 "001000110111111111101001",
						 "001000111000000001100100",
						 "001000111000000011011111",
						 "001000111000000101011010",
						 "001000111000000111010101",
						 "001000111000001001010000",
						 "001000111000001011001011",
						 "001000111000001101000110",
						 "001000111000001111000001",
						 "001000111000010000111100",
						 "001000111000010010110111",
						 "001000110111110110000010",
						 "001000110111110111111101",
						 "001000110111111001111000",
						 "001000110111111011110011",
						 "001000110111111101101110",
						 "001000110111111111101001",
						 "001000111000000001100100",
						 "001000111000000011011111",
						 "001000111000000101011010",
						 "001000111000000111010101",
						 "001000111000001001010000",
						 "001000111000001011001011",
						 "001000111000001101000110",
						 "001000111000001111000001",
						 "001000111000010000111100",
						 "001000111000010010110111",
						 "001000111010011001000000",
						 "001000111010011010111010",
						 "001000111010011100110100",
						 "001000111010011110101110",
						 "001000111010100000101000",
						 "001000111010100010100010",
						 "001000111010100100011100",
						 "001000111010100110010110",
						 "001000111010101000010000",
						 "001000111010101010001010",
						 "001000111010101100000100",
						 "001000111010101101111110",
						 "001000111010101111111000",
						 "001000111010110001110010",
						 "001000111010110011101100",
						 "001000111010110101100110",
						 "001000111010011001000000",
						 "001000111010011010111010",
						 "001000111010011100110100",
						 "001000111010011110101110",
						 "001000111010100000101000",
						 "001000111010100010100010",
						 "001000111010100100011100",
						 "001000111010100110010110",
						 "001000111010101000010000",
						 "001000111010101010001010",
						 "001000111010101100000100",
						 "001000111010101101111110",
						 "001000111010101111111000",
						 "001000111010110001110010",
						 "001000111010110011101100",
						 "001000111010110101100110",
						 "001000111010011001000000",
						 "001000111010011010111010",
						 "001000111010011100110100",
						 "001000111010011110101110",
						 "001000111010100000101000",
						 "001000111010100010100010",
						 "001000111010100100011100",
						 "001000111010100110010110",
						 "001000111010101000010000",
						 "001000111010101010001010",
						 "001000111010101100000100",
						 "001000111010101101111110",
						 "001000111010101111111000",
						 "001000111010110001110010",
						 "001000111010110011101100",
						 "001000111010110101100110",
						 "001000111010011001000000",
						 "001000111010011010111001",
						 "001000111010011100110010",
						 "001000111010011110101011",
						 "001000111010100000100100",
						 "001000111010100010011101",
						 "001000111010100100010110",
						 "001000111010100110001111",
						 "001000111010101000001000",
						 "001000111010101010000001",
						 "001000111010101011111010",
						 "001000111010101101110011",
						 "001000111010101111101100",
						 "001000111010110001100101",
						 "001000111010110011011110",
						 "001000111010110101010111",
						 "001000111010011001000000",
						 "001000111010011010111001",
						 "001000111010011100110010",
						 "001000111010011110101011",
						 "001000111010100000100100",
						 "001000111010100010011101",
						 "001000111010100100010110",
						 "001000111010100110001111",
						 "001000111010101000001000",
						 "001000111010101010000001",
						 "001000111010101011111010",
						 "001000111010101101110011",
						 "001000111010101111101100",
						 "001000111010110001100101",
						 "001000111010110011011110",
						 "001000111010110101010111",
						 "001000111100111011111110",
						 "001000111100111101110111",
						 "001000111100111111110000",
						 "001000111101000001101001",
						 "001000111101000011100010",
						 "001000111101000101011011",
						 "001000111101000111010100",
						 "001000111101001001001101",
						 "001000111101001011000110",
						 "001000111101001100111111",
						 "001000111101001110111000",
						 "001000111101010000110001",
						 "001000111101010010101010",
						 "001000111101010100100011",
						 "001000111101010110011100",
						 "001000111101011000010101",
						 "001000111100111011111110",
						 "001000111100111101110110",
						 "001000111100111111101110",
						 "001000111101000001100110",
						 "001000111101000011011110",
						 "001000111101000101010110",
						 "001000111101000111001110",
						 "001000111101001001000110",
						 "001000111101001010111110",
						 "001000111101001100110110",
						 "001000111101001110101110",
						 "001000111101010000100110",
						 "001000111101010010011110",
						 "001000111101010100010110",
						 "001000111101010110001110",
						 "001000111101011000000110",
						 "001000111100111011111110",
						 "001000111100111101110110",
						 "001000111100111111101110",
						 "001000111101000001100110",
						 "001000111101000011011110",
						 "001000111101000101010110",
						 "001000111101000111001110",
						 "001000111101001001000110",
						 "001000111101001010111110",
						 "001000111101001100110110",
						 "001000111101001110101110",
						 "001000111101010000100110",
						 "001000111101010010011110",
						 "001000111101010100010110",
						 "001000111101010110001110",
						 "001000111101011000000110",
						 "001000111100111011111110",
						 "001000111100111101110110",
						 "001000111100111111101110",
						 "001000111101000001100110",
						 "001000111101000011011110",
						 "001000111101000101010110",
						 "001000111101000111001110",
						 "001000111101001001000110",
						 "001000111101001010111110",
						 "001000111101001100110110",
						 "001000111101001110101110",
						 "001000111101010000100110",
						 "001000111101010010011110",
						 "001000111101010100010110",
						 "001000111101010110001110",
						 "001000111101011000000110",
						 "001000111100111011111110",
						 "001000111100111101110101",
						 "001000111100111111101100",
						 "001000111101000001100011",
						 "001000111101000011011010",
						 "001000111101000101010001",
						 "001000111101000111001000",
						 "001000111101001000111111",
						 "001000111101001010110110",
						 "001000111101001100101101",
						 "001000111101001110100100",
						 "001000111101010000011011",
						 "001000111101010010010010",
						 "001000111101010100001001",
						 "001000111101010110000000",
						 "001000111101010111110111",
						 "001000111100111011111110",
						 "001000111100111101110101",
						 "001000111100111111101100",
						 "001000111101000001100011",
						 "001000111101000011011010",
						 "001000111101000101010001",
						 "001000111101000111001000",
						 "001000111101001000111111",
						 "001000111101001010110110",
						 "001000111101001100101101",
						 "001000111101001110100100",
						 "001000111101010000011011",
						 "001000111101010010010010",
						 "001000111101010100001001",
						 "001000111101010110000000",
						 "001000111101010111110111",
						 "001000111111011110111100",
						 "001000111111100000110011",
						 "001000111111100010101010",
						 "001000111111100100100001",
						 "001000111111100110011000",
						 "001000111111101000001111",
						 "001000111111101010000110",
						 "001000111111101011111101",
						 "001000111111101101110100",
						 "001000111111101111101011",
						 "001000111111110001100010",
						 "001000111111110011011001",
						 "001000111111110101010000",
						 "001000111111110111000111",
						 "001000111111111000111110",
						 "001000111111111010110101",
						 "001000111111011110111100",
						 "001000111111100000110010",
						 "001000111111100010101000",
						 "001000111111100100011110",
						 "001000111111100110010100",
						 "001000111111101000001010",
						 "001000111111101010000000",
						 "001000111111101011110110",
						 "001000111111101101101100",
						 "001000111111101111100010",
						 "001000111111110001011000",
						 "001000111111110011001110",
						 "001000111111110101000100",
						 "001000111111110110111010",
						 "001000111111111000110000",
						 "001000111111111010100110",
						 "001000111111011110111100",
						 "001000111111100000110010",
						 "001000111111100010101000",
						 "001000111111100100011110",
						 "001000111111100110010100",
						 "001000111111101000001010",
						 "001000111111101010000000",
						 "001000111111101011110110",
						 "001000111111101101101100",
						 "001000111111101111100010",
						 "001000111111110001011000",
						 "001000111111110011001110",
						 "001000111111110101000100",
						 "001000111111110110111010",
						 "001000111111111000110000",
						 "001000111111111010100110",
						 "001000111111011110111100",
						 "001000111111100000110010",
						 "001000111111100010101000",
						 "001000111111100100011110",
						 "001000111111100110010100",
						 "001000111111101000001010",
						 "001000111111101010000000",
						 "001000111111101011110110",
						 "001000111111101101101100",
						 "001000111111101111100010",
						 "001000111111110001011000",
						 "001000111111110011001110",
						 "001000111111110101000100",
						 "001000111111110110111010",
						 "001000111111111000110000",
						 "001000111111111010100110",
						 "001000111111011110111100",
						 "001000111111100000110001",
						 "001000111111100010100110",
						 "001000111111100100011011",
						 "001000111111100110010000",
						 "001000111111101000000101",
						 "001000111111101001111010",
						 "001000111111101011101111",
						 "001000111111101101100100",
						 "001000111111101111011001",
						 "001000111111110001001110",
						 "001000111111110011000011",
						 "001000111111110100111000",
						 "001000111111110110101101",
						 "001000111111111000100010",
						 "001000111111111010010111",
						 "001001000010000001111010",
						 "001001000010000011101111",
						 "001001000010000101100100",
						 "001001000010000111011001",
						 "001001000010001001001110",
						 "001001000010001011000011",
						 "001001000010001100111000",
						 "001001000010001110101101",
						 "001001000010010000100010",
						 "001001000010010010010111",
						 "001001000010010100001100",
						 "001001000010010110000001",
						 "001001000010010111110110",
						 "001001000010011001101011",
						 "001001000010011011100000",
						 "001001000010011101010101",
						 "001001000010000001111010",
						 "001001000010000011101111",
						 "001001000010000101100100",
						 "001001000010000111011001",
						 "001001000010001001001110",
						 "001001000010001011000011",
						 "001001000010001100111000",
						 "001001000010001110101101",
						 "001001000010010000100010",
						 "001001000010010010010111",
						 "001001000010010100001100",
						 "001001000010010110000001",
						 "001001000010010111110110",
						 "001001000010011001101011",
						 "001001000010011011100000",
						 "001001000010011101010101",
						 "001001000010000001111010",
						 "001001000010000011101110",
						 "001001000010000101100010",
						 "001001000010000111010110",
						 "001001000010001001001010",
						 "001001000010001010111110",
						 "001001000010001100110010",
						 "001001000010001110100110",
						 "001001000010010000011010",
						 "001001000010010010001110",
						 "001001000010010100000010",
						 "001001000010010101110110",
						 "001001000010010111101010",
						 "001001000010011001011110",
						 "001001000010011011010010",
						 "001001000010011101000110",
						 "001001000010000001111010",
						 "001001000010000011101110",
						 "001001000010000101100010",
						 "001001000010000111010110",
						 "001001000010001001001010",
						 "001001000010001010111110",
						 "001001000010001100110010",
						 "001001000010001110100110",
						 "001001000010010000011010",
						 "001001000010010010001110",
						 "001001000010010100000010",
						 "001001000010010101110110",
						 "001001000010010111101010",
						 "001001000010011001011110",
						 "001001000010011011010010",
						 "001001000010011101000110",
						 "001001000010000001111010",
						 "001001000010000011101110",
						 "001001000010000101100010",
						 "001001000010000111010110",
						 "001001000010001001001010",
						 "001001000010001010111110",
						 "001001000010001100110010",
						 "001001000010001110100110",
						 "001001000010010000011010",
						 "001001000010010010001110",
						 "001001000010010100000010",
						 "001001000010010101110110",
						 "001001000010010111101010",
						 "001001000010011001011110",
						 "001001000010011011010010",
						 "001001000010011101000110",
						 "001001000010000001111010",
						 "001001000010000011101101",
						 "001001000010000101100000",
						 "001001000010000111010011",
						 "001001000010001001000110",
						 "001001000010001010111001",
						 "001001000010001100101100",
						 "001001000010001110011111",
						 "001001000010010000010010",
						 "001001000010010010000101",
						 "001001000010010011111000",
						 "001001000010010101101011",
						 "001001000010010111011110",
						 "001001000010011001010001",
						 "001001000010011011000100",
						 "001001000010011100110111",
						 "001001000100100100111000",
						 "001001000100100110101011",
						 "001001000100101000011110",
						 "001001000100101010010001",
						 "001001000100101100000100",
						 "001001000100101101110111",
						 "001001000100101111101010",
						 "001001000100110001011101",
						 "001001000100110011010000",
						 "001001000100110101000011",
						 "001001000100110110110110",
						 "001001000100111000101001",
						 "001001000100111010011100",
						 "001001000100111100001111",
						 "001001000100111110000010",
						 "001001000100111111110101",
						 "001001000100100100111000",
						 "001001000100100110101010",
						 "001001000100101000011100",
						 "001001000100101010001110",
						 "001001000100101100000000",
						 "001001000100101101110010",
						 "001001000100101111100100",
						 "001001000100110001010110",
						 "001001000100110011001000",
						 "001001000100110100111010",
						 "001001000100110110101100",
						 "001001000100111000011110",
						 "001001000100111010010000",
						 "001001000100111100000010",
						 "001001000100111101110100",
						 "001001000100111111100110",
						 "001001000100100100111000",
						 "001001000100100110101010",
						 "001001000100101000011100",
						 "001001000100101010001110",
						 "001001000100101100000000",
						 "001001000100101101110010",
						 "001001000100101111100100",
						 "001001000100110001010110",
						 "001001000100110011001000",
						 "001001000100110100111010",
						 "001001000100110110101100",
						 "001001000100111000011110",
						 "001001000100111010010000",
						 "001001000100111100000010",
						 "001001000100111101110100",
						 "001001000100111111100110",
						 "001001000100100100111000",
						 "001001000100100110101010",
						 "001001000100101000011100",
						 "001001000100101010001110",
						 "001001000100101100000000",
						 "001001000100101101110010",
						 "001001000100101111100100",
						 "001001000100110001010110",
						 "001001000100110011001000",
						 "001001000100110100111010",
						 "001001000100110110101100",
						 "001001000100111000011110",
						 "001001000100111010010000",
						 "001001000100111100000010",
						 "001001000100111101110100",
						 "001001000100111111100110",
						 "001001000100100100111000",
						 "001001000100100110101001",
						 "001001000100101000011010",
						 "001001000100101010001011",
						 "001001000100101011111100",
						 "001001000100101101101101",
						 "001001000100101111011110",
						 "001001000100110001001111",
						 "001001000100110011000000",
						 "001001000100110100110001",
						 "001001000100110110100010",
						 "001001000100111000010011",
						 "001001000100111010000100",
						 "001001000100111011110101",
						 "001001000100111101100110",
						 "001001000100111111010111",
						 "001001000100100100111000",
						 "001001000100100110101001",
						 "001001000100101000011010",
						 "001001000100101010001011",
						 "001001000100101011111100",
						 "001001000100101101101101",
						 "001001000100101111011110",
						 "001001000100110001001111",
						 "001001000100110011000000",
						 "001001000100110100110001",
						 "001001000100110110100010",
						 "001001000100111000010011",
						 "001001000100111010000100",
						 "001001000100111011110101",
						 "001001000100111101100110",
						 "001001000100111111010111",
						 "001001000111000111110110",
						 "001001000111001001100111",
						 "001001000111001011011000",
						 "001001000111001101001001",
						 "001001000111001110111010",
						 "001001000111010000101011",
						 "001001000111010010011100",
						 "001001000111010100001101",
						 "001001000111010101111110",
						 "001001000111010111101111",
						 "001001000111011001100000",
						 "001001000111011011010001",
						 "001001000111011101000010",
						 "001001000111011110110011",
						 "001001000111100000100100",
						 "001001000111100010010101",
						 "001001000111000111110110",
						 "001001000111001001100110",
						 "001001000111001011010110",
						 "001001000111001101000110",
						 "001001000111001110110110",
						 "001001000111010000100110",
						 "001001000111010010010110",
						 "001001000111010100000110",
						 "001001000111010101110110",
						 "001001000111010111100110",
						 "001001000111011001010110",
						 "001001000111011011000110",
						 "001001000111011100110110",
						 "001001000111011110100110",
						 "001001000111100000010110",
						 "001001000111100010000110",
						 "001001000111000111110110",
						 "001001000111001001100110",
						 "001001000111001011010110",
						 "001001000111001101000110",
						 "001001000111001110110110",
						 "001001000111010000100110",
						 "001001000111010010010110",
						 "001001000111010100000110",
						 "001001000111010101110110",
						 "001001000111010111100110",
						 "001001000111011001010110",
						 "001001000111011011000110",
						 "001001000111011100110110",
						 "001001000111011110100110",
						 "001001000111100000010110",
						 "001001000111100010000110",
						 "001001000111000111110110",
						 "001001000111001001100110",
						 "001001000111001011010110",
						 "001001000111001101000110",
						 "001001000111001110110110",
						 "001001000111010000100110",
						 "001001000111010010010110",
						 "001001000111010100000110",
						 "001001000111010101110110",
						 "001001000111010111100110",
						 "001001000111011001010110",
						 "001001000111011011000110",
						 "001001000111011100110110",
						 "001001000111011110100110",
						 "001001000111100000010110",
						 "001001000111100010000110",
						 "001001000111000111110110",
						 "001001000111001001100101",
						 "001001000111001011010100",
						 "001001000111001101000011",
						 "001001000111001110110010",
						 "001001000111010000100001",
						 "001001000111010010010000",
						 "001001000111010011111111",
						 "001001000111010101101110",
						 "001001000111010111011101",
						 "001001000111011001001100",
						 "001001000111011010111011",
						 "001001000111011100101010",
						 "001001000111011110011001",
						 "001001000111100000001000",
						 "001001000111100001110111",
						 "001001001001101010110100",
						 "001001001001101100100011",
						 "001001001001101110010010",
						 "001001001001110000000001",
						 "001001001001110001110000",
						 "001001001001110011011111",
						 "001001001001110101001110",
						 "001001001001110110111101",
						 "001001001001111000101100",
						 "001001001001111010011011",
						 "001001001001111100001010",
						 "001001001001111101111001",
						 "001001001001111111101000",
						 "001001001010000001010111",
						 "001001001010000011000110",
						 "001001001010000100110101",
						 "001001001001101010110100",
						 "001001001001101100100011",
						 "001001001001101110010010",
						 "001001001001110000000001",
						 "001001001001110001110000",
						 "001001001001110011011111",
						 "001001001001110101001110",
						 "001001001001110110111101",
						 "001001001001111000101100",
						 "001001001001111010011011",
						 "001001001001111100001010",
						 "001001001001111101111001",
						 "001001001001111111101000",
						 "001001001010000001010111",
						 "001001001010000011000110",
						 "001001001010000100110101",
						 "001001001001101010110100",
						 "001001001001101100100010",
						 "001001001001101110010000",
						 "001001001001101111111110",
						 "001001001001110001101100",
						 "001001001001110011011010",
						 "001001001001110101001000",
						 "001001001001110110110110",
						 "001001001001111000100100",
						 "001001001001111010010010",
						 "001001001001111100000000",
						 "001001001001111101101110",
						 "001001001001111111011100",
						 "001001001010000001001010",
						 "001001001010000010111000",
						 "001001001010000100100110",
						 "001001001001101010110100",
						 "001001001001101100100010",
						 "001001001001101110010000",
						 "001001001001101111111110",
						 "001001001001110001101100",
						 "001001001001110011011010",
						 "001001001001110101001000",
						 "001001001001110110110110",
						 "001001001001111000100100",
						 "001001001001111010010010",
						 "001001001001111100000000",
						 "001001001001111101101110",
						 "001001001001111111011100",
						 "001001001010000001001010",
						 "001001001010000010111000",
						 "001001001010000100100110",
						 "001001001001101010110100",
						 "001001001001101100100010",
						 "001001001001101110010000",
						 "001001001001101111111110",
						 "001001001001110001101100",
						 "001001001001110011011010",
						 "001001001001110101001000",
						 "001001001001110110110110",
						 "001001001001111000100100",
						 "001001001001111010010010",
						 "001001001001111100000000",
						 "001001001001111101101110",
						 "001001001001111111011100",
						 "001001001010000001001010",
						 "001001001010000010111000",
						 "001001001010000100100110",
						 "001001001001101010110100",
						 "001001001001101100100001",
						 "001001001001101110001110",
						 "001001001001101111111011",
						 "001001001001110001101000",
						 "001001001001110011010101",
						 "001001001001110101000010",
						 "001001001001110110101111",
						 "001001001001111000011100",
						 "001001001001111010001001",
						 "001001001001111011110110",
						 "001001001001111101100011",
						 "001001001001111111010000",
						 "001001001010000000111101",
						 "001001001010000010101010",
						 "001001001010000100010111",
						 "001001001100001101110010",
						 "001001001100001111011111",
						 "001001001100010001001100",
						 "001001001100010010111001",
						 "001001001100010100100110",
						 "001001001100010110010011",
						 "001001001100011000000000",
						 "001001001100011001101101",
						 "001001001100011011011010",
						 "001001001100011101000111",
						 "001001001100011110110100",
						 "001001001100100000100001",
						 "001001001100100010001110",
						 "001001001100100011111011",
						 "001001001100100101101000",
						 "001001001100100111010101",
						 "001001001100001101110010",
						 "001001001100001111011110",
						 "001001001100010001001010",
						 "001001001100010010110110",
						 "001001001100010100100010",
						 "001001001100010110001110",
						 "001001001100010111111010",
						 "001001001100011001100110",
						 "001001001100011011010010",
						 "001001001100011100111110",
						 "001001001100011110101010",
						 "001001001100100000010110",
						 "001001001100100010000010",
						 "001001001100100011101110",
						 "001001001100100101011010",
						 "001001001100100111000110",
						 "001001001100001101110010",
						 "001001001100001111011110",
						 "001001001100010001001010",
						 "001001001100010010110110",
						 "001001001100010100100010",
						 "001001001100010110001110",
						 "001001001100010111111010",
						 "001001001100011001100110",
						 "001001001100011011010010",
						 "001001001100011100111110",
						 "001001001100011110101010",
						 "001001001100100000010110",
						 "001001001100100010000010",
						 "001001001100100011101110",
						 "001001001100100101011010",
						 "001001001100100111000110",
						 "001001001100001101110010",
						 "001001001100001111011110",
						 "001001001100010001001010",
						 "001001001100010010110110",
						 "001001001100010100100010",
						 "001001001100010110001110",
						 "001001001100010111111010",
						 "001001001100011001100110",
						 "001001001100011011010010",
						 "001001001100011100111110",
						 "001001001100011110101010",
						 "001001001100100000010110",
						 "001001001100100010000010",
						 "001001001100100011101110",
						 "001001001100100101011010",
						 "001001001100100111000110",
						 "001001001100001101110010",
						 "001001001100001111011101",
						 "001001001100010001001000",
						 "001001001100010010110011",
						 "001001001100010100011110",
						 "001001001100010110001001",
						 "001001001100010111110100",
						 "001001001100011001011111",
						 "001001001100011011001010",
						 "001001001100011100110101",
						 "001001001100011110100000",
						 "001001001100100000001011",
						 "001001001100100001110110",
						 "001001001100100011100001",
						 "001001001100100101001100",
						 "001001001100100110110111",
						 "001001001100001101110010",
						 "001001001100001111011101",
						 "001001001100010001001000",
						 "001001001100010010110011",
						 "001001001100010100011110",
						 "001001001100010110001001",
						 "001001001100010111110100",
						 "001001001100011001011111",
						 "001001001100011011001010",
						 "001001001100011100110101",
						 "001001001100011110100000",
						 "001001001100100000001011",
						 "001001001100100001110110",
						 "001001001100100011100001",
						 "001001001100100101001100",
						 "001001001100100110110111",
						 "001001001110110000110000",
						 "001001001110110010011011",
						 "001001001110110100000110",
						 "001001001110110101110001",
						 "001001001110110111011100",
						 "001001001110111001000111",
						 "001001001110111010110010",
						 "001001001110111100011101",
						 "001001001110111110001000",
						 "001001001110111111110011",
						 "001001001111000001011110",
						 "001001001111000011001001",
						 "001001001111000100110100",
						 "001001001111000110011111",
						 "001001001111001000001010",
						 "001001001111001001110101",
						 "001001001110110000110000",
						 "001001001110110010011010",
						 "001001001110110100000100",
						 "001001001110110101101110",
						 "001001001110110111011000",
						 "001001001110111001000010",
						 "001001001110111010101100",
						 "001001001110111100010110",
						 "001001001110111110000000",
						 "001001001110111111101010",
						 "001001001111000001010100",
						 "001001001111000010111110",
						 "001001001111000100101000",
						 "001001001111000110010010",
						 "001001001111000111111100",
						 "001001001111001001100110",
						 "001001001110110000110000",
						 "001001001110110010011010",
						 "001001001110110100000100",
						 "001001001110110101101110",
						 "001001001110110111011000",
						 "001001001110111001000010",
						 "001001001110111010101100",
						 "001001001110111100010110",
						 "001001001110111110000000",
						 "001001001110111111101010",
						 "001001001111000001010100",
						 "001001001111000010111110",
						 "001001001111000100101000",
						 "001001001111000110010010",
						 "001001001111000111111100",
						 "001001001111001001100110",
						 "001001001110110000110000",
						 "001001001110110010011010",
						 "001001001110110100000100",
						 "001001001110110101101110",
						 "001001001110110111011000",
						 "001001001110111001000010",
						 "001001001110111010101100",
						 "001001001110111100010110",
						 "001001001110111110000000",
						 "001001001110111111101010",
						 "001001001111000001010100",
						 "001001001111000010111110",
						 "001001001111000100101000",
						 "001001001111000110010010",
						 "001001001111000111111100",
						 "001001001111001001100110",
						 "001001001110110000110000",
						 "001001001110110010011001",
						 "001001001110110100000010",
						 "001001001110110101101011",
						 "001001001110110111010100",
						 "001001001110111000111101",
						 "001001001110111010100110",
						 "001001001110111100001111",
						 "001001001110111101111000",
						 "001001001110111111100001",
						 "001001001111000001001010",
						 "001001001111000010110011",
						 "001001001111000100011100",
						 "001001001111000110000101",
						 "001001001111000111101110",
						 "001001001111001001010111",
						 "001001001110110000110000",
						 "001001001110110010011001",
						 "001001001110110100000010",
						 "001001001110110101101011",
						 "001001001110110111010100",
						 "001001001110111000111101",
						 "001001001110111010100110",
						 "001001001110111100001111",
						 "001001001110111101111000",
						 "001001001110111111100001",
						 "001001001111000001001010",
						 "001001001111000010110011",
						 "001001001111000100011100",
						 "001001001111000110000101",
						 "001001001111000111101110",
						 "001001001111001001010111",
						 "001001001110110000110000",
						 "001001001110110010011001",
						 "001001001110110100000010",
						 "001001001110110101101011",
						 "001001001110110111010100",
						 "001001001110111000111101",
						 "001001001110111010100110",
						 "001001001110111100001111",
						 "001001001110111101111000",
						 "001001001110111111100001",
						 "001001001111000001001010",
						 "001001001111000010110011",
						 "001001001111000100011100",
						 "001001001111000110000101",
						 "001001001111000111101110",
						 "001001001111001001010111",
						 "001001010001010011101110",
						 "001001010001010101010110",
						 "001001010001010110111110",
						 "001001010001011000100110",
						 "001001010001011010001110",
						 "001001010001011011110110",
						 "001001010001011101011110",
						 "001001010001011111000110",
						 "001001010001100000101110",
						 "001001010001100010010110",
						 "001001010001100011111110",
						 "001001010001100101100110",
						 "001001010001100111001110",
						 "001001010001101000110110",
						 "001001010001101010011110",
						 "001001010001101100000110",
						 "001001010001010011101110",
						 "001001010001010101010110",
						 "001001010001010110111110",
						 "001001010001011000100110",
						 "001001010001011010001110",
						 "001001010001011011110110",
						 "001001010001011101011110",
						 "001001010001011111000110",
						 "001001010001100000101110",
						 "001001010001100010010110",
						 "001001010001100011111110",
						 "001001010001100101100110",
						 "001001010001100111001110",
						 "001001010001101000110110",
						 "001001010001101010011110",
						 "001001010001101100000110",
						 "001001010001010011101110",
						 "001001010001010101010110",
						 "001001010001010110111110",
						 "001001010001011000100110",
						 "001001010001011010001110",
						 "001001010001011011110110",
						 "001001010001011101011110",
						 "001001010001011111000110",
						 "001001010001100000101110",
						 "001001010001100010010110",
						 "001001010001100011111110",
						 "001001010001100101100110",
						 "001001010001100111001110",
						 "001001010001101000110110",
						 "001001010001101010011110",
						 "001001010001101100000110",
						 "001001010001010011101110",
						 "001001010001010101010101",
						 "001001010001010110111100",
						 "001001010001011000100011",
						 "001001010001011010001010",
						 "001001010001011011110001",
						 "001001010001011101011000",
						 "001001010001011110111111",
						 "001001010001100000100110",
						 "001001010001100010001101",
						 "001001010001100011110100",
						 "001001010001100101011011",
						 "001001010001100111000010",
						 "001001010001101000101001",
						 "001001010001101010010000",
						 "001001010001101011110111",
						 "001001010001010011101110",
						 "001001010001010101010101",
						 "001001010001010110111100",
						 "001001010001011000100011",
						 "001001010001011010001010",
						 "001001010001011011110001",
						 "001001010001011101011000",
						 "001001010001011110111111",
						 "001001010001100000100110",
						 "001001010001100010001101",
						 "001001010001100011110100",
						 "001001010001100101011011",
						 "001001010001100111000010",
						 "001001010001101000101001",
						 "001001010001101010010000",
						 "001001010001101011110111",
						 "001001010001010011101110",
						 "001001010001010101010100",
						 "001001010001010110111010",
						 "001001010001011000100000",
						 "001001010001011010000110",
						 "001001010001011011101100",
						 "001001010001011101010010",
						 "001001010001011110111000",
						 "001001010001100000011110",
						 "001001010001100010000100",
						 "001001010001100011101010",
						 "001001010001100101010000",
						 "001001010001100110110110",
						 "001001010001101000011100",
						 "001001010001101010000010",
						 "001001010001101011101000",
						 "001001010011110110101100",
						 "001001010011111000010010",
						 "001001010011111001111000",
						 "001001010011111011011110",
						 "001001010011111101000100",
						 "001001010011111110101010",
						 "001001010100000000010000",
						 "001001010100000001110110",
						 "001001010100000011011100",
						 "001001010100000101000010",
						 "001001010100000110101000",
						 "001001010100001000001110",
						 "001001010100001001110100",
						 "001001010100001011011010",
						 "001001010100001101000000",
						 "001001010100001110100110",
						 "001001010011110110101100",
						 "001001010011111000010010",
						 "001001010011111001111000",
						 "001001010011111011011110",
						 "001001010011111101000100",
						 "001001010011111110101010",
						 "001001010100000000010000",
						 "001001010100000001110110",
						 "001001010100000011011100",
						 "001001010100000101000010",
						 "001001010100000110101000",
						 "001001010100001000001110",
						 "001001010100001001110100",
						 "001001010100001011011010",
						 "001001010100001101000000",
						 "001001010100001110100110",
						 "001001010011110110101100",
						 "001001010011111000010001",
						 "001001010011111001110110",
						 "001001010011111011011011",
						 "001001010011111101000000",
						 "001001010011111110100101",
						 "001001010100000000001010",
						 "001001010100000001101111",
						 "001001010100000011010100",
						 "001001010100000100111001",
						 "001001010100000110011110",
						 "001001010100001000000011",
						 "001001010100001001101000",
						 "001001010100001011001101",
						 "001001010100001100110010",
						 "001001010100001110010111",
						 "001001010011110110101100",
						 "001001010011111000010001",
						 "001001010011111001110110",
						 "001001010011111011011011",
						 "001001010011111101000000",
						 "001001010011111110100101",
						 "001001010100000000001010",
						 "001001010100000001101111",
						 "001001010100000011010100",
						 "001001010100000100111001",
						 "001001010100000110011110",
						 "001001010100001000000011",
						 "001001010100001001101000",
						 "001001010100001011001101",
						 "001001010100001100110010",
						 "001001010100001110010111",
						 "001001010011110110101100",
						 "001001010011111000010001",
						 "001001010011111001110110",
						 "001001010011111011011011",
						 "001001010011111101000000",
						 "001001010011111110100101",
						 "001001010100000000001010",
						 "001001010100000001101111",
						 "001001010100000011010100",
						 "001001010100000100111001",
						 "001001010100000110011110",
						 "001001010100001000000011",
						 "001001010100001001101000",
						 "001001010100001011001101",
						 "001001010100001100110010",
						 "001001010100001110010111",
						 "001001010011110110101100",
						 "001001010011111000010000",
						 "001001010011111001110100",
						 "001001010011111011011000",
						 "001001010011111100111100",
						 "001001010011111110100000",
						 "001001010100000000000100",
						 "001001010100000001101000",
						 "001001010100000011001100",
						 "001001010100000100110000",
						 "001001010100000110010100",
						 "001001010100000111111000",
						 "001001010100001001011100",
						 "001001010100001011000000",
						 "001001010100001100100100",
						 "001001010100001110001000",
						 "001001010110011001101010",
						 "001001010110011011001110",
						 "001001010110011100110010",
						 "001001010110011110010110",
						 "001001010110011111111010",
						 "001001010110100001011110",
						 "001001010110100011000010",
						 "001001010110100100100110",
						 "001001010110100110001010",
						 "001001010110100111101110",
						 "001001010110101001010010",
						 "001001010110101010110110",
						 "001001010110101100011010",
						 "001001010110101101111110",
						 "001001010110101111100010",
						 "001001010110110001000110",
						 "001001010110011001101010",
						 "001001010110011011001110",
						 "001001010110011100110010",
						 "001001010110011110010110",
						 "001001010110011111111010",
						 "001001010110100001011110",
						 "001001010110100011000010",
						 "001001010110100100100110",
						 "001001010110100110001010",
						 "001001010110100111101110",
						 "001001010110101001010010",
						 "001001010110101010110110",
						 "001001010110101100011010",
						 "001001010110101101111110",
						 "001001010110101111100010",
						 "001001010110110001000110",
						 "001001010110011001101010",
						 "001001010110011011001101",
						 "001001010110011100110000",
						 "001001010110011110010011",
						 "001001010110011111110110",
						 "001001010110100001011001",
						 "001001010110100010111100",
						 "001001010110100100011111",
						 "001001010110100110000010",
						 "001001010110100111100101",
						 "001001010110101001001000",
						 "001001010110101010101011",
						 "001001010110101100001110",
						 "001001010110101101110001",
						 "001001010110101111010100",
						 "001001010110110000110111",
						 "001001010110011001101010",
						 "001001010110011011001101",
						 "001001010110011100110000",
						 "001001010110011110010011",
						 "001001010110011111110110",
						 "001001010110100001011001",
						 "001001010110100010111100",
						 "001001010110100100011111",
						 "001001010110100110000010",
						 "001001010110100111100101",
						 "001001010110101001001000",
						 "001001010110101010101011",
						 "001001010110101100001110",
						 "001001010110101101110001",
						 "001001010110101111010100",
						 "001001010110110000110111",
						 "001001010110011001101010",
						 "001001010110011011001100",
						 "001001010110011100101110",
						 "001001010110011110010000",
						 "001001010110011111110010",
						 "001001010110100001010100",
						 "001001010110100010110110",
						 "001001010110100100011000",
						 "001001010110100101111010",
						 "001001010110100111011100",
						 "001001010110101000111110",
						 "001001010110101010100000",
						 "001001010110101100000010",
						 "001001010110101101100100",
						 "001001010110101111000110",
						 "001001010110110000101000",
						 "001001010110011001101010",
						 "001001010110011011001100",
						 "001001010110011100101110",
						 "001001010110011110010000",
						 "001001010110011111110010",
						 "001001010110100001010100",
						 "001001010110100010110110",
						 "001001010110100100011000",
						 "001001010110100101111010",
						 "001001010110100111011100",
						 "001001010110101000111110",
						 "001001010110101010100000",
						 "001001010110101100000010",
						 "001001010110101101100100",
						 "001001010110101111000110",
						 "001001010110110000101000",
						 "001001010110011001101010",
						 "001001010110011011001100",
						 "001001010110011100101110",
						 "001001010110011110010000",
						 "001001010110011111110010",
						 "001001010110100001010100",
						 "001001010110100010110110",
						 "001001010110100100011000",
						 "001001010110100101111010",
						 "001001010110100111011100",
						 "001001010110101000111110",
						 "001001010110101010100000",
						 "001001010110101100000010",
						 "001001010110101101100100",
						 "001001010110101111000110",
						 "001001010110110000101000",
						 "001001011000111100101000",
						 "001001011000111110001001",
						 "001001011000111111101010",
						 "001001011001000001001011",
						 "001001011001000010101100",
						 "001001011001000100001101",
						 "001001011001000101101110",
						 "001001011001000111001111",
						 "001001011001001000110000",
						 "001001011001001010010001",
						 "001001011001001011110010",
						 "001001011001001101010011",
						 "001001011001001110110100",
						 "001001011001010000010101",
						 "001001011001010001110110",
						 "001001011001010011010111",
						 "001001011000111100101000",
						 "001001011000111110001001",
						 "001001011000111111101010",
						 "001001011001000001001011",
						 "001001011001000010101100",
						 "001001011001000100001101",
						 "001001011001000101101110",
						 "001001011001000111001111",
						 "001001011001001000110000",
						 "001001011001001010010001",
						 "001001011001001011110010",
						 "001001011001001101010011",
						 "001001011001001110110100",
						 "001001011001010000010101",
						 "001001011001010001110110",
						 "001001011001010011010111",
						 "001001011000111100101000",
						 "001001011000111110001001",
						 "001001011000111111101010",
						 "001001011001000001001011",
						 "001001011001000010101100",
						 "001001011001000100001101",
						 "001001011001000101101110",
						 "001001011001000111001111",
						 "001001011001001000110000",
						 "001001011001001010010001",
						 "001001011001001011110010",
						 "001001011001001101010011",
						 "001001011001001110110100",
						 "001001011001010000010101",
						 "001001011001010001110110",
						 "001001011001010011010111",
						 "001001011000111100101000",
						 "001001011000111110001000",
						 "001001011000111111101000",
						 "001001011001000001001000",
						 "001001011001000010101000",
						 "001001011001000100001000",
						 "001001011001000101101000",
						 "001001011001000111001000",
						 "001001011001001000101000",
						 "001001011001001010001000",
						 "001001011001001011101000",
						 "001001011001001101001000",
						 "001001011001001110101000",
						 "001001011001010000001000",
						 "001001011001010001101000",
						 "001001011001010011001000",
						 "001001011000111100101000",
						 "001001011000111110001000",
						 "001001011000111111101000",
						 "001001011001000001001000",
						 "001001011001000010101000",
						 "001001011001000100001000",
						 "001001011001000101101000",
						 "001001011001000111001000",
						 "001001011001001000101000",
						 "001001011001001010001000",
						 "001001011001001011101000",
						 "001001011001001101001000",
						 "001001011001001110101000",
						 "001001011001010000001000",
						 "001001011001010001101000",
						 "001001011001010011001000",
						 "001001011000111100101000",
						 "001001011000111110001000",
						 "001001011000111111101000",
						 "001001011001000001001000",
						 "001001011001000010101000",
						 "001001011001000100001000",
						 "001001011001000101101000",
						 "001001011001000111001000",
						 "001001011001001000101000",
						 "001001011001001010001000",
						 "001001011001001011101000",
						 "001001011001001101001000",
						 "001001011001001110101000",
						 "001001011001010000001000",
						 "001001011001010001101000",
						 "001001011001010011001000",
						 "001001011000111100101000",
						 "001001011000111110000111",
						 "001001011000111111100110",
						 "001001011001000001000101",
						 "001001011001000010100100",
						 "001001011001000100000011",
						 "001001011001000101100010",
						 "001001011001000111000001",
						 "001001011001001000100000",
						 "001001011001001001111111",
						 "001001011001001011011110",
						 "001001011001001100111101",
						 "001001011001001110011100",
						 "001001011001001111111011",
						 "001001011001010001011010",
						 "001001011001010010111001",
						 "001001011011011111100110",
						 "001001011011100001000101",
						 "001001011011100010100100",
						 "001001011011100100000011",
						 "001001011011100101100010",
						 "001001011011100111000001",
						 "001001011011101000100000",
						 "001001011011101001111111",
						 "001001011011101011011110",
						 "001001011011101100111101",
						 "001001011011101110011100",
						 "001001011011101111111011",
						 "001001011011110001011010",
						 "001001011011110010111001",
						 "001001011011110100011000",
						 "001001011011110101110111",
						 "001001011011011111100110",
						 "001001011011100001000100",
						 "001001011011100010100010",
						 "001001011011100100000000",
						 "001001011011100101011110",
						 "001001011011100110111100",
						 "001001011011101000011010",
						 "001001011011101001111000",
						 "001001011011101011010110",
						 "001001011011101100110100",
						 "001001011011101110010010",
						 "001001011011101111110000",
						 "001001011011110001001110",
						 "001001011011110010101100",
						 "001001011011110100001010",
						 "001001011011110101101000",
						 "001001011011011111100110",
						 "001001011011100001000100",
						 "001001011011100010100010",
						 "001001011011100100000000",
						 "001001011011100101011110",
						 "001001011011100110111100",
						 "001001011011101000011010",
						 "001001011011101001111000",
						 "001001011011101011010110",
						 "001001011011101100110100",
						 "001001011011101110010010",
						 "001001011011101111110000",
						 "001001011011110001001110",
						 "001001011011110010101100",
						 "001001011011110100001010",
						 "001001011011110101101000",
						 "001001011011011111100110",
						 "001001011011100001000100",
						 "001001011011100010100010",
						 "001001011011100100000000",
						 "001001011011100101011110",
						 "001001011011100110111100",
						 "001001011011101000011010",
						 "001001011011101001111000",
						 "001001011011101011010110",
						 "001001011011101100110100",
						 "001001011011101110010010",
						 "001001011011101111110000",
						 "001001011011110001001110",
						 "001001011011110010101100",
						 "001001011011110100001010",
						 "001001011011110101101000",
						 "001001011011011111100110",
						 "001001011011100001000011",
						 "001001011011100010100000",
						 "001001011011100011111101",
						 "001001011011100101011010",
						 "001001011011100110110111",
						 "001001011011101000010100",
						 "001001011011101001110001",
						 "001001011011101011001110",
						 "001001011011101100101011",
						 "001001011011101110001000",
						 "001001011011101111100101",
						 "001001011011110001000010",
						 "001001011011110010011111",
						 "001001011011110011111100",
						 "001001011011110101011001",
						 "001001011011011111100110",
						 "001001011011100001000011",
						 "001001011011100010100000",
						 "001001011011100011111101",
						 "001001011011100101011010",
						 "001001011011100110110111",
						 "001001011011101000010100",
						 "001001011011101001110001",
						 "001001011011101011001110",
						 "001001011011101100101011",
						 "001001011011101110001000",
						 "001001011011101111100101",
						 "001001011011110001000010",
						 "001001011011110010011111",
						 "001001011011110011111100",
						 "001001011011110101011001",
						 "001001011011011111100110",
						 "001001011011100001000011",
						 "001001011011100010100000",
						 "001001011011100011111101",
						 "001001011011100101011010",
						 "001001011011100110110111",
						 "001001011011101000010100",
						 "001001011011101001110001",
						 "001001011011101011001110",
						 "001001011011101100101011",
						 "001001011011101110001000",
						 "001001011011101111100101",
						 "001001011011110001000010",
						 "001001011011110010011111",
						 "001001011011110011111100",
						 "001001011011110101011001",
						 "001001011110000010100100",
						 "001001011110000100000000",
						 "001001011110000101011100",
						 "001001011110000110111000",
						 "001001011110001000010100",
						 "001001011110001001110000",
						 "001001011110001011001100",
						 "001001011110001100101000",
						 "001001011110001110000100",
						 "001001011110001111100000",
						 "001001011110010000111100",
						 "001001011110010010011000",
						 "001001011110010011110100",
						 "001001011110010101010000",
						 "001001011110010110101100",
						 "001001011110011000001000",
						 "001001011110000010100100",
						 "001001011110000100000000",
						 "001001011110000101011100",
						 "001001011110000110111000",
						 "001001011110001000010100",
						 "001001011110001001110000",
						 "001001011110001011001100",
						 "001001011110001100101000",
						 "001001011110001110000100",
						 "001001011110001111100000",
						 "001001011110010000111100",
						 "001001011110010010011000",
						 "001001011110010011110100",
						 "001001011110010101010000",
						 "001001011110010110101100",
						 "001001011110011000001000",
						 "001001011110000010100100",
						 "001001011110000100000000",
						 "001001011110000101011100",
						 "001001011110000110111000",
						 "001001011110001000010100",
						 "001001011110001001110000",
						 "001001011110001011001100",
						 "001001011110001100101000",
						 "001001011110001110000100",
						 "001001011110001111100000",
						 "001001011110010000111100",
						 "001001011110010010011000",
						 "001001011110010011110100",
						 "001001011110010101010000",
						 "001001011110010110101100",
						 "001001011110011000001000",
						 "001001011110000010100100",
						 "001001011110000011111111",
						 "001001011110000101011010",
						 "001001011110000110110101",
						 "001001011110001000010000",
						 "001001011110001001101011",
						 "001001011110001011000110",
						 "001001011110001100100001",
						 "001001011110001101111100",
						 "001001011110001111010111",
						 "001001011110010000110010",
						 "001001011110010010001101",
						 "001001011110010011101000",
						 "001001011110010101000011",
						 "001001011110010110011110",
						 "001001011110010111111001",
						 "001001011110000010100100",
						 "001001011110000011111111",
						 "001001011110000101011010",
						 "001001011110000110110101",
						 "001001011110001000010000",
						 "001001011110001001101011",
						 "001001011110001011000110",
						 "001001011110001100100001",
						 "001001011110001101111100",
						 "001001011110001111010111",
						 "001001011110010000110010",
						 "001001011110010010001101",
						 "001001011110010011101000",
						 "001001011110010101000011",
						 "001001011110010110011110",
						 "001001011110010111111001",
						 "001001011110000010100100",
						 "001001011110000011111110",
						 "001001011110000101011000",
						 "001001011110000110110010",
						 "001001011110001000001100",
						 "001001011110001001100110",
						 "001001011110001011000000",
						 "001001011110001100011010",
						 "001001011110001101110100",
						 "001001011110001111001110",
						 "001001011110010000101000",
						 "001001011110010010000010",
						 "001001011110010011011100",
						 "001001011110010100110110",
						 "001001011110010110010000",
						 "001001011110010111101010",
						 "001001011110000010100100",
						 "001001011110000011111110",
						 "001001011110000101011000",
						 "001001011110000110110010",
						 "001001011110001000001100",
						 "001001011110001001100110",
						 "001001011110001011000000",
						 "001001011110001100011010",
						 "001001011110001101110100",
						 "001001011110001111001110",
						 "001001011110010000101000",
						 "001001011110010010000010",
						 "001001011110010011011100",
						 "001001011110010100110110",
						 "001001011110010110010000",
						 "001001011110010111101010",
						 "001001100000100101100010",
						 "001001100000100110111100",
						 "001001100000101000010110",
						 "001001100000101001110000",
						 "001001100000101011001010",
						 "001001100000101100100100",
						 "001001100000101101111110",
						 "001001100000101111011000",
						 "001001100000110000110010",
						 "001001100000110010001100",
						 "001001100000110011100110",
						 "001001100000110101000000",
						 "001001100000110110011010",
						 "001001100000110111110100",
						 "001001100000111001001110",
						 "001001100000111010101000",
						 "001001100000100101100010",
						 "001001100000100110111011",
						 "001001100000101000010100",
						 "001001100000101001101101",
						 "001001100000101011000110",
						 "001001100000101100011111",
						 "001001100000101101111000",
						 "001001100000101111010001",
						 "001001100000110000101010",
						 "001001100000110010000011",
						 "001001100000110011011100",
						 "001001100000110100110101",
						 "001001100000110110001110",
						 "001001100000110111100111",
						 "001001100000111001000000",
						 "001001100000111010011001",
						 "001001100000100101100010",
						 "001001100000100110111011",
						 "001001100000101000010100",
						 "001001100000101001101101",
						 "001001100000101011000110",
						 "001001100000101100011111",
						 "001001100000101101111000",
						 "001001100000101111010001",
						 "001001100000110000101010",
						 "001001100000110010000011",
						 "001001100000110011011100",
						 "001001100000110100110101",
						 "001001100000110110001110",
						 "001001100000110111100111",
						 "001001100000111001000000",
						 "001001100000111010011001",
						 "001001100000100101100010",
						 "001001100000100110111011",
						 "001001100000101000010100",
						 "001001100000101001101101",
						 "001001100000101011000110",
						 "001001100000101100011111",
						 "001001100000101101111000",
						 "001001100000101111010001",
						 "001001100000110000101010",
						 "001001100000110010000011",
						 "001001100000110011011100",
						 "001001100000110100110101",
						 "001001100000110110001110",
						 "001001100000110111100111",
						 "001001100000111001000000",
						 "001001100000111010011001",
						 "001001100000100101100010",
						 "001001100000100110111010",
						 "001001100000101000010010",
						 "001001100000101001101010",
						 "001001100000101011000010",
						 "001001100000101100011010",
						 "001001100000101101110010",
						 "001001100000101111001010",
						 "001001100000110000100010",
						 "001001100000110001111010",
						 "001001100000110011010010",
						 "001001100000110100101010",
						 "001001100000110110000010",
						 "001001100000110111011010",
						 "001001100000111000110010",
						 "001001100000111010001010",
						 "001001100000100101100010",
						 "001001100000100110111010",
						 "001001100000101000010010",
						 "001001100000101001101010",
						 "001001100000101011000010",
						 "001001100000101100011010",
						 "001001100000101101110010",
						 "001001100000101111001010",
						 "001001100000110000100010",
						 "001001100000110001111010",
						 "001001100000110011010010",
						 "001001100000110100101010",
						 "001001100000110110000010",
						 "001001100000110111011010",
						 "001001100000111000110010",
						 "001001100000111010001010",
						 "001001100000100101100010",
						 "001001100000100110111010",
						 "001001100000101000010010",
						 "001001100000101001101010",
						 "001001100000101011000010",
						 "001001100000101100011010",
						 "001001100000101101110010",
						 "001001100000101111001010",
						 "001001100000110000100010",
						 "001001100000110001111010",
						 "001001100000110011010010",
						 "001001100000110100101010",
						 "001001100000110110000010",
						 "001001100000110111011010",
						 "001001100000111000110010",
						 "001001100000111010001010",
						 "001001100011001000100000",
						 "001001100011001001110111",
						 "001001100011001011001110",
						 "001001100011001100100101",
						 "001001100011001101111100",
						 "001001100011001111010011",
						 "001001100011010000101010",
						 "001001100011010010000001",
						 "001001100011010011011000",
						 "001001100011010100101111",
						 "001001100011010110000110",
						 "001001100011010111011101",
						 "001001100011011000110100",
						 "001001100011011010001011",
						 "001001100011011011100010",
						 "001001100011011100111001",
						 "001001100011001000100000",
						 "001001100011001001110111",
						 "001001100011001011001110",
						 "001001100011001100100101",
						 "001001100011001101111100",
						 "001001100011001111010011",
						 "001001100011010000101010",
						 "001001100011010010000001",
						 "001001100011010011011000",
						 "001001100011010100101111",
						 "001001100011010110000110",
						 "001001100011010111011101",
						 "001001100011011000110100",
						 "001001100011011010001011",
						 "001001100011011011100010",
						 "001001100011011100111001",
						 "001001100011001000100000",
						 "001001100011001001110110",
						 "001001100011001011001100",
						 "001001100011001100100010",
						 "001001100011001101111000",
						 "001001100011001111001110",
						 "001001100011010000100100",
						 "001001100011010001111010",
						 "001001100011010011010000",
						 "001001100011010100100110",
						 "001001100011010101111100",
						 "001001100011010111010010",
						 "001001100011011000101000",
						 "001001100011011001111110",
						 "001001100011011011010100",
						 "001001100011011100101010",
						 "001001100011001000100000",
						 "001001100011001001110110",
						 "001001100011001011001100",
						 "001001100011001100100010",
						 "001001100011001101111000",
						 "001001100011001111001110",
						 "001001100011010000100100",
						 "001001100011010001111010",
						 "001001100011010011010000",
						 "001001100011010100100110",
						 "001001100011010101111100",
						 "001001100011010111010010",
						 "001001100011011000101000",
						 "001001100011011001111110",
						 "001001100011011011010100",
						 "001001100011011100101010",
						 "001001100011001000100000",
						 "001001100011001001110110",
						 "001001100011001011001100",
						 "001001100011001100100010",
						 "001001100011001101111000",
						 "001001100011001111001110",
						 "001001100011010000100100",
						 "001001100011010001111010",
						 "001001100011010011010000",
						 "001001100011010100100110",
						 "001001100011010101111100",
						 "001001100011010111010010",
						 "001001100011011000101000",
						 "001001100011011001111110",
						 "001001100011011011010100",
						 "001001100011011100101010",
						 "001001100011001000100000",
						 "001001100011001001110101",
						 "001001100011001011001010",
						 "001001100011001100011111",
						 "001001100011001101110100",
						 "001001100011001111001001",
						 "001001100011010000011110",
						 "001001100011010001110011",
						 "001001100011010011001000",
						 "001001100011010100011101",
						 "001001100011010101110010",
						 "001001100011010111000111",
						 "001001100011011000011100",
						 "001001100011011001110001",
						 "001001100011011011000110",
						 "001001100011011100011011",
						 "001001100011001000100000",
						 "001001100011001001110101",
						 "001001100011001011001010",
						 "001001100011001100011111",
						 "001001100011001101110100",
						 "001001100011001111001001",
						 "001001100011010000011110",
						 "001001100011010001110011",
						 "001001100011010011001000",
						 "001001100011010100011101",
						 "001001100011010101110010",
						 "001001100011010111000111",
						 "001001100011011000011100",
						 "001001100011011001110001",
						 "001001100011011011000110",
						 "001001100011011100011011",
						 "001001100011001000100000",
						 "001001100011001001110101",
						 "001001100011001011001010",
						 "001001100011001100011111",
						 "001001100011001101110100",
						 "001001100011001111001001",
						 "001001100011010000011110",
						 "001001100011010001110011",
						 "001001100011010011001000",
						 "001001100011010100011101",
						 "001001100011010101110010",
						 "001001100011010111000111",
						 "001001100011011000011100",
						 "001001100011011001110001",
						 "001001100011011011000110",
						 "001001100011011100011011",
						 "001001100101101011011110",
						 "001001100101101100110010",
						 "001001100101101110000110",
						 "001001100101101111011010",
						 "001001100101110000101110",
						 "001001100101110010000010",
						 "001001100101110011010110",
						 "001001100101110100101010",
						 "001001100101110101111110",
						 "001001100101110111010010",
						 "001001100101111000100110",
						 "001001100101111001111010",
						 "001001100101111011001110",
						 "001001100101111100100010",
						 "001001100101111101110110",
						 "001001100101111111001010",
						 "001001100101101011011110",
						 "001001100101101100110010",
						 "001001100101101110000110",
						 "001001100101101111011010",
						 "001001100101110000101110",
						 "001001100101110010000010",
						 "001001100101110011010110",
						 "001001100101110100101010",
						 "001001100101110101111110",
						 "001001100101110111010010",
						 "001001100101111000100110",
						 "001001100101111001111010",
						 "001001100101111011001110",
						 "001001100101111100100010",
						 "001001100101111101110110",
						 "001001100101111111001010",
						 "001001100101101011011110",
						 "001001100101101100110001",
						 "001001100101101110000100",
						 "001001100101101111010111",
						 "001001100101110000101010",
						 "001001100101110001111101",
						 "001001100101110011010000",
						 "001001100101110100100011",
						 "001001100101110101110110",
						 "001001100101110111001001",
						 "001001100101111000011100",
						 "001001100101111001101111",
						 "001001100101111011000010",
						 "001001100101111100010101",
						 "001001100101111101101000",
						 "001001100101111110111011",
						 "001001100101101011011110",
						 "001001100101101100110001",
						 "001001100101101110000100",
						 "001001100101101111010111",
						 "001001100101110000101010",
						 "001001100101110001111101",
						 "001001100101110011010000",
						 "001001100101110100100011",
						 "001001100101110101110110",
						 "001001100101110111001001",
						 "001001100101111000011100",
						 "001001100101111001101111",
						 "001001100101111011000010",
						 "001001100101111100010101",
						 "001001100101111101101000",
						 "001001100101111110111011",
						 "001001100101101011011110",
						 "001001100101101100110001",
						 "001001100101101110000100",
						 "001001100101101111010111",
						 "001001100101110000101010",
						 "001001100101110001111101",
						 "001001100101110011010000",
						 "001001100101110100100011",
						 "001001100101110101110110",
						 "001001100101110111001001",
						 "001001100101111000011100",
						 "001001100101111001101111",
						 "001001100101111011000010",
						 "001001100101111100010101",
						 "001001100101111101101000",
						 "001001100101111110111011",
						 "001001100101101011011110",
						 "001001100101101100110000",
						 "001001100101101110000010",
						 "001001100101101111010100",
						 "001001100101110000100110",
						 "001001100101110001111000",
						 "001001100101110011001010",
						 "001001100101110100011100",
						 "001001100101110101101110",
						 "001001100101110111000000",
						 "001001100101111000010010",
						 "001001100101111001100100",
						 "001001100101111010110110",
						 "001001100101111100001000",
						 "001001100101111101011010",
						 "001001100101111110101100",
						 "001001100101101011011110",
						 "001001100101101100110000",
						 "001001100101101110000010",
						 "001001100101101111010100",
						 "001001100101110000100110",
						 "001001100101110001111000",
						 "001001100101110011001010",
						 "001001100101110100011100",
						 "001001100101110101101110",
						 "001001100101110111000000",
						 "001001100101111000010010",
						 "001001100101111001100100",
						 "001001100101111010110110",
						 "001001100101111100001000",
						 "001001100101111101011010",
						 "001001100101111110101100",
						 "001001101000001110011100",
						 "001001101000001111101110",
						 "001001101000010001000000",
						 "001001101000010010010010",
						 "001001101000010011100100",
						 "001001101000010100110110",
						 "001001101000010110001000",
						 "001001101000010111011010",
						 "001001101000011000101100",
						 "001001101000011001111110",
						 "001001101000011011010000",
						 "001001101000011100100010",
						 "001001101000011101110100",
						 "001001101000011111000110",
						 "001001101000100000011000",
						 "001001101000100001101010",
						 "001001101000001110011100",
						 "001001101000001111101101",
						 "001001101000010000111110",
						 "001001101000010010001111",
						 "001001101000010011100000",
						 "001001101000010100110001",
						 "001001101000010110000010",
						 "001001101000010111010011",
						 "001001101000011000100100",
						 "001001101000011001110101",
						 "001001101000011011000110",
						 "001001101000011100010111",
						 "001001101000011101101000",
						 "001001101000011110111001",
						 "001001101000100000001010",
						 "001001101000100001011011",
						 "001001101000001110011100",
						 "001001101000001111101101",
						 "001001101000010000111110",
						 "001001101000010010001111",
						 "001001101000010011100000",
						 "001001101000010100110001",
						 "001001101000010110000010",
						 "001001101000010111010011",
						 "001001101000011000100100",
						 "001001101000011001110101",
						 "001001101000011011000110",
						 "001001101000011100010111",
						 "001001101000011101101000",
						 "001001101000011110111001",
						 "001001101000100000001010",
						 "001001101000100001011011",
						 "001001101000001110011100",
						 "001001101000001111101101",
						 "001001101000010000111110",
						 "001001101000010010001111",
						 "001001101000010011100000",
						 "001001101000010100110001",
						 "001001101000010110000010",
						 "001001101000010111010011",
						 "001001101000011000100100",
						 "001001101000011001110101",
						 "001001101000011011000110",
						 "001001101000011100010111",
						 "001001101000011101101000",
						 "001001101000011110111001",
						 "001001101000100000001010",
						 "001001101000100001011011",
						 "001001101000001110011100",
						 "001001101000001111101100",
						 "001001101000010000111100",
						 "001001101000010010001100",
						 "001001101000010011011100",
						 "001001101000010100101100",
						 "001001101000010101111100",
						 "001001101000010111001100",
						 "001001101000011000011100",
						 "001001101000011001101100",
						 "001001101000011010111100",
						 "001001101000011100001100",
						 "001001101000011101011100",
						 "001001101000011110101100",
						 "001001101000011111111100",
						 "001001101000100001001100",
						 "001001101000001110011100",
						 "001001101000001111101100",
						 "001001101000010000111100",
						 "001001101000010010001100",
						 "001001101000010011011100",
						 "001001101000010100101100",
						 "001001101000010101111100",
						 "001001101000010111001100",
						 "001001101000011000011100",
						 "001001101000011001101100",
						 "001001101000011010111100",
						 "001001101000011100001100",
						 "001001101000011101011100",
						 "001001101000011110101100",
						 "001001101000011111111100",
						 "001001101000100001001100",
						 "001001101000001110011100",
						 "001001101000001111101011",
						 "001001101000010000111010",
						 "001001101000010010001001",
						 "001001101000010011011000",
						 "001001101000010100100111",
						 "001001101000010101110110",
						 "001001101000010111000101",
						 "001001101000011000010100",
						 "001001101000011001100011",
						 "001001101000011010110010",
						 "001001101000011100000001",
						 "001001101000011101010000",
						 "001001101000011110011111",
						 "001001101000011111101110",
						 "001001101000100000111101",
						 "001001101000001110011100",
						 "001001101000001111101011",
						 "001001101000010000111010",
						 "001001101000010010001001",
						 "001001101000010011011000",
						 "001001101000010100100111",
						 "001001101000010101110110",
						 "001001101000010111000101",
						 "001001101000011000010100",
						 "001001101000011001100011",
						 "001001101000011010110010",
						 "001001101000011100000001",
						 "001001101000011101010000",
						 "001001101000011110011111",
						 "001001101000011111101110",
						 "001001101000100000111101",
						 "001001101000001110011100",
						 "001001101000001111101011",
						 "001001101000010000111010",
						 "001001101000010010001001",
						 "001001101000010011011000",
						 "001001101000010100100111",
						 "001001101000010101110110",
						 "001001101000010111000101",
						 "001001101000011000010100",
						 "001001101000011001100011",
						 "001001101000011010110010",
						 "001001101000011100000001",
						 "001001101000011101010000",
						 "001001101000011110011111",
						 "001001101000011111101110",
						 "001001101000100000111101",
						 "001001101010110001011010",
						 "001001101010110010101000",
						 "001001101010110011110110",
						 "001001101010110101000100",
						 "001001101010110110010010",
						 "001001101010110111100000",
						 "001001101010111000101110",
						 "001001101010111001111100",
						 "001001101010111011001010",
						 "001001101010111100011000",
						 "001001101010111101100110",
						 "001001101010111110110100",
						 "001001101011000000000010",
						 "001001101011000001010000",
						 "001001101011000010011110",
						 "001001101011000011101100",
						 "001001101010110001011010",
						 "001001101010110010101000",
						 "001001101010110011110110",
						 "001001101010110101000100",
						 "001001101010110110010010",
						 "001001101010110111100000",
						 "001001101010111000101110",
						 "001001101010111001111100",
						 "001001101010111011001010",
						 "001001101010111100011000",
						 "001001101010111101100110",
						 "001001101010111110110100",
						 "001001101011000000000010",
						 "001001101011000001010000",
						 "001001101011000010011110",
						 "001001101011000011101100",
						 "001001101010110001011010",
						 "001001101010110010101000",
						 "001001101010110011110110",
						 "001001101010110101000100",
						 "001001101010110110010010",
						 "001001101010110111100000",
						 "001001101010111000101110",
						 "001001101010111001111100",
						 "001001101010111011001010",
						 "001001101010111100011000",
						 "001001101010111101100110",
						 "001001101010111110110100",
						 "001001101011000000000010",
						 "001001101011000001010000",
						 "001001101011000010011110",
						 "001001101011000011101100",
						 "001001101010110001011010",
						 "001001101010110010100111",
						 "001001101010110011110100",
						 "001001101010110101000001",
						 "001001101010110110001110",
						 "001001101010110111011011",
						 "001001101010111000101000",
						 "001001101010111001110101",
						 "001001101010111011000010",
						 "001001101010111100001111",
						 "001001101010111101011100",
						 "001001101010111110101001",
						 "001001101010111111110110",
						 "001001101011000001000011",
						 "001001101011000010010000",
						 "001001101011000011011101",
						 "001001101010110001011010",
						 "001001101010110010100111",
						 "001001101010110011110100",
						 "001001101010110101000001",
						 "001001101010110110001110",
						 "001001101010110111011011",
						 "001001101010111000101000",
						 "001001101010111001110101",
						 "001001101010111011000010",
						 "001001101010111100001111",
						 "001001101010111101011100",
						 "001001101010111110101001",
						 "001001101010111111110110",
						 "001001101011000001000011",
						 "001001101011000010010000",
						 "001001101011000011011101",
						 "001001101010110001011010",
						 "001001101010110010100110",
						 "001001101010110011110010",
						 "001001101010110100111110",
						 "001001101010110110001010",
						 "001001101010110111010110",
						 "001001101010111000100010",
						 "001001101010111001101110",
						 "001001101010111010111010",
						 "001001101010111100000110",
						 "001001101010111101010010",
						 "001001101010111110011110",
						 "001001101010111111101010",
						 "001001101011000000110110",
						 "001001101011000010000010",
						 "001001101011000011001110",
						 "001001101010110001011010",
						 "001001101010110010100110",
						 "001001101010110011110010",
						 "001001101010110100111110",
						 "001001101010110110001010",
						 "001001101010110111010110",
						 "001001101010111000100010",
						 "001001101010111001101110",
						 "001001101010111010111010",
						 "001001101010111100000110",
						 "001001101010111101010010",
						 "001001101010111110011110",
						 "001001101010111111101010",
						 "001001101011000000110110",
						 "001001101011000010000010",
						 "001001101011000011001110",
						 "001001101010110001011010",
						 "001001101010110010100110",
						 "001001101010110011110010",
						 "001001101010110100111110",
						 "001001101010110110001010",
						 "001001101010110111010110",
						 "001001101010111000100010",
						 "001001101010111001101110",
						 "001001101010111010111010",
						 "001001101010111100000110",
						 "001001101010111101010010",
						 "001001101010111110011110",
						 "001001101010111111101010",
						 "001001101011000000110110",
						 "001001101011000010000010",
						 "001001101011000011001110",
						 "001001101101010100011000",
						 "001001101101010101100011",
						 "001001101101010110101110",
						 "001001101101010111111001",
						 "001001101101011001000100",
						 "001001101101011010001111",
						 "001001101101011011011010",
						 "001001101101011100100101",
						 "001001101101011101110000",
						 "001001101101011110111011",
						 "001001101101100000000110",
						 "001001101101100001010001",
						 "001001101101100010011100",
						 "001001101101100011100111",
						 "001001101101100100110010",
						 "001001101101100101111101",
						 "001001101101010100011000",
						 "001001101101010101100011",
						 "001001101101010110101110",
						 "001001101101010111111001",
						 "001001101101011001000100",
						 "001001101101011010001111",
						 "001001101101011011011010",
						 "001001101101011100100101",
						 "001001101101011101110000",
						 "001001101101011110111011",
						 "001001101101100000000110",
						 "001001101101100001010001",
						 "001001101101100010011100",
						 "001001101101100011100111",
						 "001001101101100100110010",
						 "001001101101100101111101",
						 "001001101101010100011000",
						 "001001101101010101100011",
						 "001001101101010110101110",
						 "001001101101010111111001",
						 "001001101101011001000100",
						 "001001101101011010001111",
						 "001001101101011011011010",
						 "001001101101011100100101",
						 "001001101101011101110000",
						 "001001101101011110111011",
						 "001001101101100000000110",
						 "001001101101100001010001",
						 "001001101101100010011100",
						 "001001101101100011100111",
						 "001001101101100100110010",
						 "001001101101100101111101",
						 "001001101101010100011000",
						 "001001101101010101100010",
						 "001001101101010110101100",
						 "001001101101010111110110",
						 "001001101101011001000000",
						 "001001101101011010001010",
						 "001001101101011011010100",
						 "001001101101011100011110",
						 "001001101101011101101000",
						 "001001101101011110110010",
						 "001001101101011111111100",
						 "001001101101100001000110",
						 "001001101101100010010000",
						 "001001101101100011011010",
						 "001001101101100100100100",
						 "001001101101100101101110",
						 "001001101101010100011000",
						 "001001101101010101100010",
						 "001001101101010110101100",
						 "001001101101010111110110",
						 "001001101101011001000000",
						 "001001101101011010001010",
						 "001001101101011011010100",
						 "001001101101011100011110",
						 "001001101101011101101000",
						 "001001101101011110110010",
						 "001001101101011111111100",
						 "001001101101100001000110",
						 "001001101101100010010000",
						 "001001101101100011011010",
						 "001001101101100100100100",
						 "001001101101100101101110",
						 "001001101101010100011000",
						 "001001101101010101100001",
						 "001001101101010110101010",
						 "001001101101010111110011",
						 "001001101101011000111100",
						 "001001101101011010000101",
						 "001001101101011011001110",
						 "001001101101011100010111",
						 "001001101101011101100000",
						 "001001101101011110101001",
						 "001001101101011111110010",
						 "001001101101100000111011",
						 "001001101101100010000100",
						 "001001101101100011001101",
						 "001001101101100100010110",
						 "001001101101100101011111",
						 "001001101101010100011000",
						 "001001101101010101100001",
						 "001001101101010110101010",
						 "001001101101010111110011",
						 "001001101101011000111100",
						 "001001101101011010000101",
						 "001001101101011011001110",
						 "001001101101011100010111",
						 "001001101101011101100000",
						 "001001101101011110101001",
						 "001001101101011111110010",
						 "001001101101100000111011",
						 "001001101101100010000100",
						 "001001101101100011001101",
						 "001001101101100100010110",
						 "001001101101100101011111",
						 "001001101101010100011000",
						 "001001101101010101100001",
						 "001001101101010110101010",
						 "001001101101010111110011",
						 "001001101101011000111100",
						 "001001101101011010000101",
						 "001001101101011011001110",
						 "001001101101011100010111",
						 "001001101101011101100000",
						 "001001101101011110101001",
						 "001001101101011111110010",
						 "001001101101100000111011",
						 "001001101101100010000100",
						 "001001101101100011001101",
						 "001001101101100100010110",
						 "001001101101100101011111",
						 "001001101101010100011000",
						 "001001101101010101100000",
						 "001001101101010110101000",
						 "001001101101010111110000",
						 "001001101101011000111000",
						 "001001101101011010000000",
						 "001001101101011011001000",
						 "001001101101011100010000",
						 "001001101101011101011000",
						 "001001101101011110100000",
						 "001001101101011111101000",
						 "001001101101100000110000",
						 "001001101101100001111000",
						 "001001101101100011000000",
						 "001001101101100100001000",
						 "001001101101100101010000",
						 "001001101111110111010110",
						 "001001101111111000011110",
						 "001001101111111001100110",
						 "001001101111111010101110",
						 "001001101111111011110110",
						 "001001101111111100111110",
						 "001001101111111110000110",
						 "001001101111111111001110",
						 "001001110000000000010110",
						 "001001110000000001011110",
						 "001001110000000010100110",
						 "001001110000000011101110",
						 "001001110000000100110110",
						 "001001110000000101111110",
						 "001001110000000111000110",
						 "001001110000001000001110",
						 "001001101111110111010110",
						 "001001101111111000011110",
						 "001001101111111001100110",
						 "001001101111111010101110",
						 "001001101111111011110110",
						 "001001101111111100111110",
						 "001001101111111110000110",
						 "001001101111111111001110",
						 "001001110000000000010110",
						 "001001110000000001011110",
						 "001001110000000010100110",
						 "001001110000000011101110",
						 "001001110000000100110110",
						 "001001110000000101111110",
						 "001001110000000111000110",
						 "001001110000001000001110",
						 "001001101111110111010110",
						 "001001101111111000011101",
						 "001001101111111001100100",
						 "001001101111111010101011",
						 "001001101111111011110010",
						 "001001101111111100111001",
						 "001001101111111110000000",
						 "001001101111111111000111",
						 "001001110000000000001110",
						 "001001110000000001010101",
						 "001001110000000010011100",
						 "001001110000000011100011",
						 "001001110000000100101010",
						 "001001110000000101110001",
						 "001001110000000110111000",
						 "001001110000000111111111",
						 "001001101111110111010110",
						 "001001101111111000011101",
						 "001001101111111001100100",
						 "001001101111111010101011",
						 "001001101111111011110010",
						 "001001101111111100111001",
						 "001001101111111110000000",
						 "001001101111111111000111",
						 "001001110000000000001110",
						 "001001110000000001010101",
						 "001001110000000010011100",
						 "001001110000000011100011",
						 "001001110000000100101010",
						 "001001110000000101110001",
						 "001001110000000110111000",
						 "001001110000000111111111",
						 "001001101111110111010110",
						 "001001101111111000011100",
						 "001001101111111001100010",
						 "001001101111111010101000",
						 "001001101111111011101110",
						 "001001101111111100110100",
						 "001001101111111101111010",
						 "001001101111111111000000",
						 "001001110000000000000110",
						 "001001110000000001001100",
						 "001001110000000010010010",
						 "001001110000000011011000",
						 "001001110000000100011110",
						 "001001110000000101100100",
						 "001001110000000110101010",
						 "001001110000000111110000",
						 "001001101111110111010110",
						 "001001101111111000011100",
						 "001001101111111001100010",
						 "001001101111111010101000",
						 "001001101111111011101110",
						 "001001101111111100110100",
						 "001001101111111101111010",
						 "001001101111111111000000",
						 "001001110000000000000110",
						 "001001110000000001001100",
						 "001001110000000010010010",
						 "001001110000000011011000",
						 "001001110000000100011110",
						 "001001110000000101100100",
						 "001001110000000110101010",
						 "001001110000000111110000",
						 "001001101111110111010110",
						 "001001101111111000011100",
						 "001001101111111001100010",
						 "001001101111111010101000",
						 "001001101111111011101110",
						 "001001101111111100110100",
						 "001001101111111101111010",
						 "001001101111111111000000",
						 "001001110000000000000110",
						 "001001110000000001001100",
						 "001001110000000010010010",
						 "001001110000000011011000",
						 "001001110000000100011110",
						 "001001110000000101100100",
						 "001001110000000110101010",
						 "001001110000000111110000",
						 "001001101111110111010110",
						 "001001101111111000011011",
						 "001001101111111001100000",
						 "001001101111111010100101",
						 "001001101111111011101010",
						 "001001101111111100101111",
						 "001001101111111101110100",
						 "001001101111111110111001",
						 "001001101111111111111110",
						 "001001110000000001000011",
						 "001001110000000010001000",
						 "001001110000000011001101",
						 "001001110000000100010010",
						 "001001110000000101010111",
						 "001001110000000110011100",
						 "001001110000000111100001",
						 "001001101111110111010110",
						 "001001101111111000011011",
						 "001001101111111001100000",
						 "001001101111111010100101",
						 "001001101111111011101010",
						 "001001101111111100101111",
						 "001001101111111101110100",
						 "001001101111111110111001",
						 "001001101111111111111110",
						 "001001110000000001000011",
						 "001001110000000010001000",
						 "001001110000000011001101",
						 "001001110000000100010010",
						 "001001110000000101010111",
						 "001001110000000110011100",
						 "001001110000000111100001",
						 "001001110010011010010100",
						 "001001110010011011011001",
						 "001001110010011100011110",
						 "001001110010011101100011",
						 "001001110010011110101000",
						 "001001110010011111101101",
						 "001001110010100000110010",
						 "001001110010100001110111",
						 "001001110010100010111100",
						 "001001110010100100000001",
						 "001001110010100101000110",
						 "001001110010100110001011",
						 "001001110010100111010000",
						 "001001110010101000010101",
						 "001001110010101001011010",
						 "001001110010101010011111",
						 "001001110010011010010100",
						 "001001110010011011011000",
						 "001001110010011100011100",
						 "001001110010011101100000",
						 "001001110010011110100100",
						 "001001110010011111101000",
						 "001001110010100000101100",
						 "001001110010100001110000",
						 "001001110010100010110100",
						 "001001110010100011111000",
						 "001001110010100100111100",
						 "001001110010100110000000",
						 "001001110010100111000100",
						 "001001110010101000001000",
						 "001001110010101001001100",
						 "001001110010101010010000",
						 "001001110010011010010100",
						 "001001110010011011011000",
						 "001001110010011100011100",
						 "001001110010011101100000",
						 "001001110010011110100100",
						 "001001110010011111101000",
						 "001001110010100000101100",
						 "001001110010100001110000",
						 "001001110010100010110100",
						 "001001110010100011111000",
						 "001001110010100100111100",
						 "001001110010100110000000",
						 "001001110010100111000100",
						 "001001110010101000001000",
						 "001001110010101001001100",
						 "001001110010101010010000",
						 "001001110010011010010100",
						 "001001110010011011010111",
						 "001001110010011100011010",
						 "001001110010011101011101",
						 "001001110010011110100000",
						 "001001110010011111100011",
						 "001001110010100000100110",
						 "001001110010100001101001",
						 "001001110010100010101100",
						 "001001110010100011101111",
						 "001001110010100100110010",
						 "001001110010100101110101",
						 "001001110010100110111000",
						 "001001110010100111111011",
						 "001001110010101000111110",
						 "001001110010101010000001",
						 "001001110010011010010100",
						 "001001110010011011010111",
						 "001001110010011100011010",
						 "001001110010011101011101",
						 "001001110010011110100000",
						 "001001110010011111100011",
						 "001001110010100000100110",
						 "001001110010100001101001",
						 "001001110010100010101100",
						 "001001110010100011101111",
						 "001001110010100100110010",
						 "001001110010100101110101",
						 "001001110010100110111000",
						 "001001110010100111111011",
						 "001001110010101000111110",
						 "001001110010101010000001",
						 "001001110010011010010100",
						 "001001110010011011010111",
						 "001001110010011100011010",
						 "001001110010011101011101",
						 "001001110010011110100000",
						 "001001110010011111100011",
						 "001001110010100000100110",
						 "001001110010100001101001",
						 "001001110010100010101100",
						 "001001110010100011101111",
						 "001001110010100100110010",
						 "001001110010100101110101",
						 "001001110010100110111000",
						 "001001110010100111111011",
						 "001001110010101000111110",
						 "001001110010101010000001",
						 "001001110010011010010100",
						 "001001110010011011010110",
						 "001001110010011100011000",
						 "001001110010011101011010",
						 "001001110010011110011100",
						 "001001110010011111011110",
						 "001001110010100000100000",
						 "001001110010100001100010",
						 "001001110010100010100100",
						 "001001110010100011100110",
						 "001001110010100100101000",
						 "001001110010100101101010",
						 "001001110010100110101100",
						 "001001110010100111101110",
						 "001001110010101000110000",
						 "001001110010101001110010",
						 "001001110010011010010100",
						 "001001110010011011010110",
						 "001001110010011100011000",
						 "001001110010011101011010",
						 "001001110010011110011100",
						 "001001110010011111011110",
						 "001001110010100000100000",
						 "001001110010100001100010",
						 "001001110010100010100100",
						 "001001110010100011100110",
						 "001001110010100100101000",
						 "001001110010100101101010",
						 "001001110010100110101100",
						 "001001110010100111101110",
						 "001001110010101000110000",
						 "001001110010101001110010",
						 "001001110010011010010100",
						 "001001110010011011010110",
						 "001001110010011100011000",
						 "001001110010011101011010",
						 "001001110010011110011100",
						 "001001110010011111011110",
						 "001001110010100000100000",
						 "001001110010100001100010",
						 "001001110010100010100100",
						 "001001110010100011100110",
						 "001001110010100100101000",
						 "001001110010100101101010",
						 "001001110010100110101100",
						 "001001110010100111101110",
						 "001001110010101000110000",
						 "001001110010101001110010",
						 "001001110010011010010100",
						 "001001110010011011010101",
						 "001001110010011100010110",
						 "001001110010011101010111",
						 "001001110010011110011000",
						 "001001110010011111011001",
						 "001001110010100000011010",
						 "001001110010100001011011",
						 "001001110010100010011100",
						 "001001110010100011011101",
						 "001001110010100100011110",
						 "001001110010100101011111",
						 "001001110010100110100000",
						 "001001110010100111100001",
						 "001001110010101000100010",
						 "001001110010101001100011",
						 "001001110100111101010010",
						 "001001110100111110010011",
						 "001001110100111111010100",
						 "001001110101000000010101",
						 "001001110101000001010110",
						 "001001110101000010010111",
						 "001001110101000011011000",
						 "001001110101000100011001",
						 "001001110101000101011010",
						 "001001110101000110011011",
						 "001001110101000111011100",
						 "001001110101001000011101",
						 "001001110101001001011110",
						 "001001110101001010011111",
						 "001001110101001011100000",
						 "001001110101001100100001",
						 "001001110100111101010010",
						 "001001110100111110010010",
						 "001001110100111111010010",
						 "001001110101000000010010",
						 "001001110101000001010010",
						 "001001110101000010010010",
						 "001001110101000011010010",
						 "001001110101000100010010",
						 "001001110101000101010010",
						 "001001110101000110010010",
						 "001001110101000111010010",
						 "001001110101001000010010",
						 "001001110101001001010010",
						 "001001110101001010010010",
						 "001001110101001011010010",
						 "001001110101001100010010",
						 "001001110100111101010010",
						 "001001110100111110010010",
						 "001001110100111111010010",
						 "001001110101000000010010",
						 "001001110101000001010010",
						 "001001110101000010010010",
						 "001001110101000011010010",
						 "001001110101000100010010",
						 "001001110101000101010010",
						 "001001110101000110010010",
						 "001001110101000111010010",
						 "001001110101001000010010",
						 "001001110101001001010010",
						 "001001110101001010010010",
						 "001001110101001011010010",
						 "001001110101001100010010",
						 "001001110100111101010010",
						 "001001110100111110010010",
						 "001001110100111111010010",
						 "001001110101000000010010",
						 "001001110101000001010010",
						 "001001110101000010010010",
						 "001001110101000011010010",
						 "001001110101000100010010",
						 "001001110101000101010010",
						 "001001110101000110010010",
						 "001001110101000111010010",
						 "001001110101001000010010",
						 "001001110101001001010010",
						 "001001110101001010010010",
						 "001001110101001011010010",
						 "001001110101001100010010",
						 "001001110100111101010010",
						 "001001110100111110010001",
						 "001001110100111111010000",
						 "001001110101000000001111",
						 "001001110101000001001110",
						 "001001110101000010001101",
						 "001001110101000011001100",
						 "001001110101000100001011",
						 "001001110101000101001010",
						 "001001110101000110001001",
						 "001001110101000111001000",
						 "001001110101001000000111",
						 "001001110101001001000110",
						 "001001110101001010000101",
						 "001001110101001011000100",
						 "001001110101001100000011",
						 "001001110100111101010010",
						 "001001110100111110010001",
						 "001001110100111111010000",
						 "001001110101000000001111",
						 "001001110101000001001110",
						 "001001110101000010001101",
						 "001001110101000011001100",
						 "001001110101000100001011",
						 "001001110101000101001010",
						 "001001110101000110001001",
						 "001001110101000111001000",
						 "001001110101001000000111",
						 "001001110101001001000110",
						 "001001110101001010000101",
						 "001001110101001011000100",
						 "001001110101001100000011",
						 "001001110100111101010010",
						 "001001110100111110010001",
						 "001001110100111111010000",
						 "001001110101000000001111",
						 "001001110101000001001110",
						 "001001110101000010001101",
						 "001001110101000011001100",
						 "001001110101000100001011",
						 "001001110101000101001010",
						 "001001110101000110001001",
						 "001001110101000111001000",
						 "001001110101001000000111",
						 "001001110101001001000110",
						 "001001110101001010000101",
						 "001001110101001011000100",
						 "001001110101001100000011",
						 "001001110100111101010010",
						 "001001110100111110010000",
						 "001001110100111111001110",
						 "001001110101000000001100",
						 "001001110101000001001010",
						 "001001110101000010001000",
						 "001001110101000011000110",
						 "001001110101000100000100",
						 "001001110101000101000010",
						 "001001110101000110000000",
						 "001001110101000110111110",
						 "001001110101000111111100",
						 "001001110101001000111010",
						 "001001110101001001111000",
						 "001001110101001010110110",
						 "001001110101001011110100",
						 "001001110100111101010010",
						 "001001110100111110010000",
						 "001001110100111111001110",
						 "001001110101000000001100",
						 "001001110101000001001010",
						 "001001110101000010001000",
						 "001001110101000011000110",
						 "001001110101000100000100",
						 "001001110101000101000010",
						 "001001110101000110000000",
						 "001001110101000110111110",
						 "001001110101000111111100",
						 "001001110101001000111010",
						 "001001110101001001111000",
						 "001001110101001010110110",
						 "001001110101001011110100",
						 "001001110100111101010010",
						 "001001110100111110001111",
						 "001001110100111111001100",
						 "001001110101000000001001",
						 "001001110101000001000110",
						 "001001110101000010000011",
						 "001001110101000011000000",
						 "001001110101000011111101",
						 "001001110101000100111010",
						 "001001110101000101110111",
						 "001001110101000110110100",
						 "001001110101000111110001",
						 "001001110101001000101110",
						 "001001110101001001101011",
						 "001001110101001010101000",
						 "001001110101001011100101",
						 "001001110111100000010000",
						 "001001110111100001001101",
						 "001001110111100010001010",
						 "001001110111100011000111",
						 "001001110111100100000100",
						 "001001110111100101000001",
						 "001001110111100101111110",
						 "001001110111100110111011",
						 "001001110111100111111000",
						 "001001110111101000110101",
						 "001001110111101001110010",
						 "001001110111101010101111",
						 "001001110111101011101100",
						 "001001110111101100101001",
						 "001001110111101101100110",
						 "001001110111101110100011",
						 "001001110111100000010000",
						 "001001110111100001001101",
						 "001001110111100010001010",
						 "001001110111100011000111",
						 "001001110111100100000100",
						 "001001110111100101000001",
						 "001001110111100101111110",
						 "001001110111100110111011",
						 "001001110111100111111000",
						 "001001110111101000110101",
						 "001001110111101001110010",
						 "001001110111101010101111",
						 "001001110111101011101100",
						 "001001110111101100101001",
						 "001001110111101101100110",
						 "001001110111101110100011",
						 "001001110111100000010000",
						 "001001110111100001001100",
						 "001001110111100010001000",
						 "001001110111100011000100",
						 "001001110111100100000000",
						 "001001110111100100111100",
						 "001001110111100101111000",
						 "001001110111100110110100",
						 "001001110111100111110000",
						 "001001110111101000101100",
						 "001001110111101001101000",
						 "001001110111101010100100",
						 "001001110111101011100000",
						 "001001110111101100011100",
						 "001001110111101101011000",
						 "001001110111101110010100",
						 "001001110111100000010000",
						 "001001110111100001001100",
						 "001001110111100010001000",
						 "001001110111100011000100",
						 "001001110111100100000000",
						 "001001110111100100111100",
						 "001001110111100101111000",
						 "001001110111100110110100",
						 "001001110111100111110000",
						 "001001110111101000101100",
						 "001001110111101001101000",
						 "001001110111101010100100",
						 "001001110111101011100000",
						 "001001110111101100011100",
						 "001001110111101101011000",
						 "001001110111101110010100",
						 "001001110111100000010000",
						 "001001110111100001001011",
						 "001001110111100010000110",
						 "001001110111100011000001",
						 "001001110111100011111100",
						 "001001110111100100110111",
						 "001001110111100101110010",
						 "001001110111100110101101",
						 "001001110111100111101000",
						 "001001110111101000100011",
						 "001001110111101001011110",
						 "001001110111101010011001",
						 "001001110111101011010100",
						 "001001110111101100001111",
						 "001001110111101101001010",
						 "001001110111101110000101",
						 "001001110111100000010000",
						 "001001110111100001001011",
						 "001001110111100010000110",
						 "001001110111100011000001",
						 "001001110111100011111100",
						 "001001110111100100110111",
						 "001001110111100101110010",
						 "001001110111100110101101",
						 "001001110111100111101000",
						 "001001110111101000100011",
						 "001001110111101001011110",
						 "001001110111101010011001",
						 "001001110111101011010100",
						 "001001110111101100001111",
						 "001001110111101101001010",
						 "001001110111101110000101",
						 "001001110111100000010000",
						 "001001110111100001001011",
						 "001001110111100010000110",
						 "001001110111100011000001",
						 "001001110111100011111100",
						 "001001110111100100110111",
						 "001001110111100101110010",
						 "001001110111100110101101",
						 "001001110111100111101000",
						 "001001110111101000100011",
						 "001001110111101001011110",
						 "001001110111101010011001",
						 "001001110111101011010100",
						 "001001110111101100001111",
						 "001001110111101101001010",
						 "001001110111101110000101",
						 "001001110111100000010000",
						 "001001110111100001001010",
						 "001001110111100010000100",
						 "001001110111100010111110",
						 "001001110111100011111000",
						 "001001110111100100110010",
						 "001001110111100101101100",
						 "001001110111100110100110",
						 "001001110111100111100000",
						 "001001110111101000011010",
						 "001001110111101001010100",
						 "001001110111101010001110",
						 "001001110111101011001000",
						 "001001110111101100000010",
						 "001001110111101100111100",
						 "001001110111101101110110",
						 "001001110111100000010000",
						 "001001110111100001001010",
						 "001001110111100010000100",
						 "001001110111100010111110",
						 "001001110111100011111000",
						 "001001110111100100110010",
						 "001001110111100101101100",
						 "001001110111100110100110",
						 "001001110111100111100000",
						 "001001110111101000011010",
						 "001001110111101001010100",
						 "001001110111101010001110",
						 "001001110111101011001000",
						 "001001110111101100000010",
						 "001001110111101100111100",
						 "001001110111101101110110",
						 "001001110111100000010000",
						 "001001110111100001001010",
						 "001001110111100010000100",
						 "001001110111100010111110",
						 "001001110111100011111000",
						 "001001110111100100110010",
						 "001001110111100101101100",
						 "001001110111100110100110",
						 "001001110111100111100000",
						 "001001110111101000011010",
						 "001001110111101001010100",
						 "001001110111101010001110",
						 "001001110111101011001000",
						 "001001110111101100000010",
						 "001001110111101100111100",
						 "001001110111101101110110",
						 "001001110111100000010000",
						 "001001110111100001001001",
						 "001001110111100010000010",
						 "001001110111100010111011",
						 "001001110111100011110100",
						 "001001110111100100101101",
						 "001001110111100101100110",
						 "001001110111100110011111",
						 "001001110111100111011000",
						 "001001110111101000010001",
						 "001001110111101001001010",
						 "001001110111101010000011",
						 "001001110111101010111100",
						 "001001110111101011110101",
						 "001001110111101100101110",
						 "001001110111101101100111",
						 "001001111010000011001110",
						 "001001111010000100000111",
						 "001001111010000101000000",
						 "001001111010000101111001",
						 "001001111010000110110010",
						 "001001111010000111101011",
						 "001001111010001000100100",
						 "001001111010001001011101",
						 "001001111010001010010110",
						 "001001111010001011001111",
						 "001001111010001100001000",
						 "001001111010001101000001",
						 "001001111010001101111010",
						 "001001111010001110110011",
						 "001001111010001111101100",
						 "001001111010010000100101",
						 "001001111010000011001110",
						 "001001111010000100000110",
						 "001001111010000100111110",
						 "001001111010000101110110",
						 "001001111010000110101110",
						 "001001111010000111100110",
						 "001001111010001000011110",
						 "001001111010001001010110",
						 "001001111010001010001110",
						 "001001111010001011000110",
						 "001001111010001011111110",
						 "001001111010001100110110",
						 "001001111010001101101110",
						 "001001111010001110100110",
						 "001001111010001111011110",
						 "001001111010010000010110",
						 "001001111010000011001110",
						 "001001111010000100000110",
						 "001001111010000100111110",
						 "001001111010000101110110",
						 "001001111010000110101110",
						 "001001111010000111100110",
						 "001001111010001000011110",
						 "001001111010001001010110",
						 "001001111010001010001110",
						 "001001111010001011000110",
						 "001001111010001011111110",
						 "001001111010001100110110",
						 "001001111010001101101110",
						 "001001111010001110100110",
						 "001001111010001111011110",
						 "001001111010010000010110",
						 "001001111010000011001110",
						 "001001111010000100000110",
						 "001001111010000100111110",
						 "001001111010000101110110",
						 "001001111010000110101110",
						 "001001111010000111100110",
						 "001001111010001000011110",
						 "001001111010001001010110",
						 "001001111010001010001110",
						 "001001111010001011000110",
						 "001001111010001011111110",
						 "001001111010001100110110",
						 "001001111010001101101110",
						 "001001111010001110100110",
						 "001001111010001111011110",
						 "001001111010010000010110",
						 "001001111010000011001110",
						 "001001111010000100000101",
						 "001001111010000100111100",
						 "001001111010000101110011",
						 "001001111010000110101010",
						 "001001111010000111100001",
						 "001001111010001000011000",
						 "001001111010001001001111",
						 "001001111010001010000110",
						 "001001111010001010111101",
						 "001001111010001011110100",
						 "001001111010001100101011",
						 "001001111010001101100010",
						 "001001111010001110011001",
						 "001001111010001111010000",
						 "001001111010010000000111",
						 "001001111010000011001110",
						 "001001111010000100000101",
						 "001001111010000100111100",
						 "001001111010000101110011",
						 "001001111010000110101010",
						 "001001111010000111100001",
						 "001001111010001000011000",
						 "001001111010001001001111",
						 "001001111010001010000110",
						 "001001111010001010111101",
						 "001001111010001011110100",
						 "001001111010001100101011",
						 "001001111010001101100010",
						 "001001111010001110011001",
						 "001001111010001111010000",
						 "001001111010010000000111",
						 "001001111010000011001110",
						 "001001111010000100000101",
						 "001001111010000100111100",
						 "001001111010000101110011",
						 "001001111010000110101010",
						 "001001111010000111100001",
						 "001001111010001000011000",
						 "001001111010001001001111",
						 "001001111010001010000110",
						 "001001111010001010111101",
						 "001001111010001011110100",
						 "001001111010001100101011",
						 "001001111010001101100010",
						 "001001111010001110011001",
						 "001001111010001111010000",
						 "001001111010010000000111",
						 "001001111010000011001110",
						 "001001111010000100000100",
						 "001001111010000100111010",
						 "001001111010000101110000",
						 "001001111010000110100110",
						 "001001111010000111011100",
						 "001001111010001000010010",
						 "001001111010001001001000",
						 "001001111010001001111110",
						 "001001111010001010110100",
						 "001001111010001011101010",
						 "001001111010001100100000",
						 "001001111010001101010110",
						 "001001111010001110001100",
						 "001001111010001111000010",
						 "001001111010001111111000",
						 "001001111010000011001110",
						 "001001111010000100000100",
						 "001001111010000100111010",
						 "001001111010000101110000",
						 "001001111010000110100110",
						 "001001111010000111011100",
						 "001001111010001000010010",
						 "001001111010001001001000",
						 "001001111010001001111110",
						 "001001111010001010110100",
						 "001001111010001011101010",
						 "001001111010001100100000",
						 "001001111010001101010110",
						 "001001111010001110001100",
						 "001001111010001111000010",
						 "001001111010001111111000",
						 "001001111010000011001110",
						 "001001111010000100000011",
						 "001001111010000100111000",
						 "001001111010000101101101",
						 "001001111010000110100010",
						 "001001111010000111010111",
						 "001001111010001000001100",
						 "001001111010001001000001",
						 "001001111010001001110110",
						 "001001111010001010101011",
						 "001001111010001011100000",
						 "001001111010001100010101",
						 "001001111010001101001010",
						 "001001111010001101111111",
						 "001001111010001110110100",
						 "001001111010001111101001",
						 "001001111010000011001110",
						 "001001111010000100000011",
						 "001001111010000100111000",
						 "001001111010000101101101",
						 "001001111010000110100010",
						 "001001111010000111010111",
						 "001001111010001000001100",
						 "001001111010001001000001",
						 "001001111010001001110110",
						 "001001111010001010101011",
						 "001001111010001011100000",
						 "001001111010001100010101",
						 "001001111010001101001010",
						 "001001111010001101111111",
						 "001001111010001110110100",
						 "001001111010001111101001",
						 "001001111010000011001110",
						 "001001111010000100000011",
						 "001001111010000100111000",
						 "001001111010000101101101",
						 "001001111010000110100010",
						 "001001111010000111010111",
						 "001001111010001000001100",
						 "001001111010001001000001",
						 "001001111010001001110110",
						 "001001111010001010101011",
						 "001001111010001011100000",
						 "001001111010001100010101",
						 "001001111010001101001010",
						 "001001111010001101111111",
						 "001001111010001110110100",
						 "001001111010001111101001",
						 "001001111100100110001100",
						 "001001111100100111000000",
						 "001001111100100111110100",
						 "001001111100101000101000",
						 "001001111100101001011100",
						 "001001111100101010010000",
						 "001001111100101011000100",
						 "001001111100101011111000",
						 "001001111100101100101100",
						 "001001111100101101100000",
						 "001001111100101110010100",
						 "001001111100101111001000",
						 "001001111100101111111100",
						 "001001111100110000110000",
						 "001001111100110001100100",
						 "001001111100110010011000",
						 "001001111100100110001100",
						 "001001111100100111000000",
						 "001001111100100111110100",
						 "001001111100101000101000",
						 "001001111100101001011100",
						 "001001111100101010010000",
						 "001001111100101011000100",
						 "001001111100101011111000",
						 "001001111100101100101100",
						 "001001111100101101100000",
						 "001001111100101110010100",
						 "001001111100101111001000",
						 "001001111100101111111100",
						 "001001111100110000110000",
						 "001001111100110001100100",
						 "001001111100110010011000",
						 "001001111100100110001100",
						 "001001111100100110111111",
						 "001001111100100111110010",
						 "001001111100101000100101",
						 "001001111100101001011000",
						 "001001111100101010001011",
						 "001001111100101010111110",
						 "001001111100101011110001",
						 "001001111100101100100100",
						 "001001111100101101010111",
						 "001001111100101110001010",
						 "001001111100101110111101",
						 "001001111100101111110000",
						 "001001111100110000100011",
						 "001001111100110001010110",
						 "001001111100110010001001",
						 "001001111100100110001100",
						 "001001111100100110111111",
						 "001001111100100111110010",
						 "001001111100101000100101",
						 "001001111100101001011000",
						 "001001111100101010001011",
						 "001001111100101010111110",
						 "001001111100101011110001",
						 "001001111100101100100100",
						 "001001111100101101010111",
						 "001001111100101110001010",
						 "001001111100101110111101",
						 "001001111100101111110000",
						 "001001111100110000100011",
						 "001001111100110001010110",
						 "001001111100110010001001",
						 "001001111100100110001100",
						 "001001111100100110111111",
						 "001001111100100111110010",
						 "001001111100101000100101",
						 "001001111100101001011000",
						 "001001111100101010001011",
						 "001001111100101010111110",
						 "001001111100101011110001",
						 "001001111100101100100100",
						 "001001111100101101010111",
						 "001001111100101110001010",
						 "001001111100101110111101",
						 "001001111100101111110000",
						 "001001111100110000100011",
						 "001001111100110001010110",
						 "001001111100110010001001",
						 "001001111100100110001100",
						 "001001111100100110111110",
						 "001001111100100111110000",
						 "001001111100101000100010",
						 "001001111100101001010100",
						 "001001111100101010000110",
						 "001001111100101010111000",
						 "001001111100101011101010",
						 "001001111100101100011100",
						 "001001111100101101001110",
						 "001001111100101110000000",
						 "001001111100101110110010",
						 "001001111100101111100100",
						 "001001111100110000010110",
						 "001001111100110001001000",
						 "001001111100110001111010",
						 "001001111100100110001100",
						 "001001111100100110111110",
						 "001001111100100111110000",
						 "001001111100101000100010",
						 "001001111100101001010100",
						 "001001111100101010000110",
						 "001001111100101010111000",
						 "001001111100101011101010",
						 "001001111100101100011100",
						 "001001111100101101001110",
						 "001001111100101110000000",
						 "001001111100101110110010",
						 "001001111100101111100100",
						 "001001111100110000010110",
						 "001001111100110001001000",
						 "001001111100110001111010",
						 "001001111100100110001100",
						 "001001111100100110111110",
						 "001001111100100111110000",
						 "001001111100101000100010",
						 "001001111100101001010100",
						 "001001111100101010000110",
						 "001001111100101010111000",
						 "001001111100101011101010",
						 "001001111100101100011100",
						 "001001111100101101001110",
						 "001001111100101110000000",
						 "001001111100101110110010",
						 "001001111100101111100100",
						 "001001111100110000010110",
						 "001001111100110001001000",
						 "001001111100110001111010",
						 "001001111100100110001100",
						 "001001111100100110111101",
						 "001001111100100111101110",
						 "001001111100101000011111",
						 "001001111100101001010000",
						 "001001111100101010000001",
						 "001001111100101010110010",
						 "001001111100101011100011",
						 "001001111100101100010100",
						 "001001111100101101000101",
						 "001001111100101101110110",
						 "001001111100101110100111",
						 "001001111100101111011000",
						 "001001111100110000001001",
						 "001001111100110000111010",
						 "001001111100110001101011",
						 "001001111100100110001100",
						 "001001111100100110111101",
						 "001001111100100111101110",
						 "001001111100101000011111",
						 "001001111100101001010000",
						 "001001111100101010000001",
						 "001001111100101010110010",
						 "001001111100101011100011",
						 "001001111100101100010100",
						 "001001111100101101000101",
						 "001001111100101101110110",
						 "001001111100101110100111",
						 "001001111100101111011000",
						 "001001111100110000001001",
						 "001001111100110000111010",
						 "001001111100110001101011",
						 "001001111100100110001100",
						 "001001111100100110111100",
						 "001001111100100111101100",
						 "001001111100101000011100",
						 "001001111100101001001100",
						 "001001111100101001111100",
						 "001001111100101010101100",
						 "001001111100101011011100",
						 "001001111100101100001100",
						 "001001111100101100111100",
						 "001001111100101101101100",
						 "001001111100101110011100",
						 "001001111100101111001100",
						 "001001111100101111111100",
						 "001001111100110000101100",
						 "001001111100110001011100",
						 "001001111100100110001100",
						 "001001111100100110111100",
						 "001001111100100111101100",
						 "001001111100101000011100",
						 "001001111100101001001100",
						 "001001111100101001111100",
						 "001001111100101010101100",
						 "001001111100101011011100",
						 "001001111100101100001100",
						 "001001111100101100111100",
						 "001001111100101101101100",
						 "001001111100101110011100",
						 "001001111100101111001100",
						 "001001111100101111111100",
						 "001001111100110000101100",
						 "001001111100110001011100",
						 "001001111100100110001100",
						 "001001111100100110111100",
						 "001001111100100111101100",
						 "001001111100101000011100",
						 "001001111100101001001100",
						 "001001111100101001111100",
						 "001001111100101010101100",
						 "001001111100101011011100",
						 "001001111100101100001100",
						 "001001111100101100111100",
						 "001001111100101101101100",
						 "001001111100101110011100",
						 "001001111100101111001100",
						 "001001111100101111111100",
						 "001001111100110000101100",
						 "001001111100110001011100",
						 "001001111111001001001010",
						 "001001111111001001111001",
						 "001001111111001010101000",
						 "001001111111001011010111",
						 "001001111111001100000110",
						 "001001111111001100110101",
						 "001001111111001101100100",
						 "001001111111001110010011",
						 "001001111111001111000010",
						 "001001111111001111110001",
						 "001001111111010000100000",
						 "001001111111010001001111",
						 "001001111111010001111110",
						 "001001111111010010101101",
						 "001001111111010011011100",
						 "001001111111010100001011",
						 "001001111111001001001010",
						 "001001111111001001111001",
						 "001001111111001010101000",
						 "001001111111001011010111",
						 "001001111111001100000110",
						 "001001111111001100110101",
						 "001001111111001101100100",
						 "001001111111001110010011",
						 "001001111111001111000010",
						 "001001111111001111110001",
						 "001001111111010000100000",
						 "001001111111010001001111",
						 "001001111111010001111110",
						 "001001111111010010101101",
						 "001001111111010011011100",
						 "001001111111010100001011",
						 "001001111111001001001010",
						 "001001111111001001111000",
						 "001001111111001010100110",
						 "001001111111001011010100",
						 "001001111111001100000010",
						 "001001111111001100110000",
						 "001001111111001101011110",
						 "001001111111001110001100",
						 "001001111111001110111010",
						 "001001111111001111101000",
						 "001001111111010000010110",
						 "001001111111010001000100",
						 "001001111111010001110010",
						 "001001111111010010100000",
						 "001001111111010011001110",
						 "001001111111010011111100",
						 "001001111111001001001010",
						 "001001111111001001111000",
						 "001001111111001010100110",
						 "001001111111001011010100",
						 "001001111111001100000010",
						 "001001111111001100110000",
						 "001001111111001101011110",
						 "001001111111001110001100",
						 "001001111111001110111010",
						 "001001111111001111101000",
						 "001001111111010000010110",
						 "001001111111010001000100",
						 "001001111111010001110010",
						 "001001111111010010100000",
						 "001001111111010011001110",
						 "001001111111010011111100",
						 "001001111111001001001010",
						 "001001111111001001111000",
						 "001001111111001010100110",
						 "001001111111001011010100",
						 "001001111111001100000010",
						 "001001111111001100110000",
						 "001001111111001101011110",
						 "001001111111001110001100",
						 "001001111111001110111010",
						 "001001111111001111101000",
						 "001001111111010000010110",
						 "001001111111010001000100",
						 "001001111111010001110010",
						 "001001111111010010100000",
						 "001001111111010011001110",
						 "001001111111010011111100",
						 "001001111111001001001010",
						 "001001111111001001110111",
						 "001001111111001010100100",
						 "001001111111001011010001",
						 "001001111111001011111110",
						 "001001111111001100101011",
						 "001001111111001101011000",
						 "001001111111001110000101",
						 "001001111111001110110010",
						 "001001111111001111011111",
						 "001001111111010000001100",
						 "001001111111010000111001",
						 "001001111111010001100110",
						 "001001111111010010010011",
						 "001001111111010011000000",
						 "001001111111010011101101",
						 "001001111111001001001010",
						 "001001111111001001110111",
						 "001001111111001010100100",
						 "001001111111001011010001",
						 "001001111111001011111110",
						 "001001111111001100101011",
						 "001001111111001101011000",
						 "001001111111001110000101",
						 "001001111111001110110010",
						 "001001111111001111011111",
						 "001001111111010000001100",
						 "001001111111010000111001",
						 "001001111111010001100110",
						 "001001111111010010010011",
						 "001001111111010011000000",
						 "001001111111010011101101",
						 "001001111111001001001010",
						 "001001111111001001110111",
						 "001001111111001010100100",
						 "001001111111001011010001",
						 "001001111111001011111110",
						 "001001111111001100101011",
						 "001001111111001101011000",
						 "001001111111001110000101",
						 "001001111111001110110010",
						 "001001111111001111011111",
						 "001001111111010000001100",
						 "001001111111010000111001",
						 "001001111111010001100110",
						 "001001111111010010010011",
						 "001001111111010011000000",
						 "001001111111010011101101",
						 "001001111111001001001010",
						 "001001111111001001110110",
						 "001001111111001010100010",
						 "001001111111001011001110",
						 "001001111111001011111010",
						 "001001111111001100100110",
						 "001001111111001101010010",
						 "001001111111001101111110",
						 "001001111111001110101010",
						 "001001111111001111010110",
						 "001001111111010000000010",
						 "001001111111010000101110",
						 "001001111111010001011010",
						 "001001111111010010000110",
						 "001001111111010010110010",
						 "001001111111010011011110",
						 "001001111111001001001010",
						 "001001111111001001110110",
						 "001001111111001010100010",
						 "001001111111001011001110",
						 "001001111111001011111010",
						 "001001111111001100100110",
						 "001001111111001101010010",
						 "001001111111001101111110",
						 "001001111111001110101010",
						 "001001111111001111010110",
						 "001001111111010000000010",
						 "001001111111010000101110",
						 "001001111111010001011010",
						 "001001111111010010000110",
						 "001001111111010010110010",
						 "001001111111010011011110",
						 "001001111111001001001010",
						 "001001111111001001110101",
						 "001001111111001010100000",
						 "001001111111001011001011",
						 "001001111111001011110110",
						 "001001111111001100100001",
						 "001001111111001101001100",
						 "001001111111001101110111",
						 "001001111111001110100010",
						 "001001111111001111001101",
						 "001001111111001111111000",
						 "001001111111010000100011",
						 "001001111111010001001110",
						 "001001111111010001111001",
						 "001001111111010010100100",
						 "001001111111010011001111",
						 "001001111111001001001010",
						 "001001111111001001110101",
						 "001001111111001010100000",
						 "001001111111001011001011",
						 "001001111111001011110110",
						 "001001111111001100100001",
						 "001001111111001101001100",
						 "001001111111001101110111",
						 "001001111111001110100010",
						 "001001111111001111001101",
						 "001001111111001111111000",
						 "001001111111010000100011",
						 "001001111111010001001110",
						 "001001111111010001111001",
						 "001001111111010010100100",
						 "001001111111010011001111",
						 "001001111111001001001010",
						 "001001111111001001110101",
						 "001001111111001010100000",
						 "001001111111001011001011",
						 "001001111111001011110110",
						 "001001111111001100100001",
						 "001001111111001101001100",
						 "001001111111001101110111",
						 "001001111111001110100010",
						 "001001111111001111001101",
						 "001001111111001111111000",
						 "001001111111010000100011",
						 "001001111111010001001110",
						 "001001111111010001111001",
						 "001001111111010010100100",
						 "001001111111010011001111",
						 "001001111111001001001010",
						 "001001111111001001110100",
						 "001001111111001010011110",
						 "001001111111001011001000",
						 "001001111111001011110010",
						 "001001111111001100011100",
						 "001001111111001101000110",
						 "001001111111001101110000",
						 "001001111111001110011010",
						 "001001111111001111000100",
						 "001001111111001111101110",
						 "001001111111010000011000",
						 "001001111111010001000010",
						 "001001111111010001101100",
						 "001001111111010010010110",
						 "001001111111010011000000",
						 "001010000001101100001000",
						 "001010000001101100110010",
						 "001010000001101101011100",
						 "001010000001101110000110",
						 "001010000001101110110000",
						 "001010000001101111011010",
						 "001010000001110000000100",
						 "001010000001110000101110",
						 "001010000001110001011000",
						 "001010000001110010000010",
						 "001010000001110010101100",
						 "001010000001110011010110",
						 "001010000001110100000000",
						 "001010000001110100101010",
						 "001010000001110101010100",
						 "001010000001110101111110",
						 "001010000001101100001000",
						 "001010000001101100110001",
						 "001010000001101101011010",
						 "001010000001101110000011",
						 "001010000001101110101100",
						 "001010000001101111010101",
						 "001010000001101111111110",
						 "001010000001110000100111",
						 "001010000001110001010000",
						 "001010000001110001111001",
						 "001010000001110010100010",
						 "001010000001110011001011",
						 "001010000001110011110100",
						 "001010000001110100011101",
						 "001010000001110101000110",
						 "001010000001110101101111",
						 "001010000001101100001000",
						 "001010000001101100110001",
						 "001010000001101101011010",
						 "001010000001101110000011",
						 "001010000001101110101100",
						 "001010000001101111010101",
						 "001010000001101111111110",
						 "001010000001110000100111",
						 "001010000001110001010000",
						 "001010000001110001111001",
						 "001010000001110010100010",
						 "001010000001110011001011",
						 "001010000001110011110100",
						 "001010000001110100011101",
						 "001010000001110101000110",
						 "001010000001110101101111",
						 "001010000001101100001000",
						 "001010000001101100110001",
						 "001010000001101101011010",
						 "001010000001101110000011",
						 "001010000001101110101100",
						 "001010000001101111010101",
						 "001010000001101111111110",
						 "001010000001110000100111",
						 "001010000001110001010000",
						 "001010000001110001111001",
						 "001010000001110010100010",
						 "001010000001110011001011",
						 "001010000001110011110100",
						 "001010000001110100011101",
						 "001010000001110101000110",
						 "001010000001110101101111",
						 "001010000001101100001000",
						 "001010000001101100110000",
						 "001010000001101101011000",
						 "001010000001101110000000",
						 "001010000001101110101000",
						 "001010000001101111010000",
						 "001010000001101111111000",
						 "001010000001110000100000",
						 "001010000001110001001000",
						 "001010000001110001110000",
						 "001010000001110010011000",
						 "001010000001110011000000",
						 "001010000001110011101000",
						 "001010000001110100010000",
						 "001010000001110100111000",
						 "001010000001110101100000",
						 "001010000001101100001000",
						 "001010000001101100110000",
						 "001010000001101101011000",
						 "001010000001101110000000",
						 "001010000001101110101000",
						 "001010000001101111010000",
						 "001010000001101111111000",
						 "001010000001110000100000",
						 "001010000001110001001000",
						 "001010000001110001110000",
						 "001010000001110010011000",
						 "001010000001110011000000",
						 "001010000001110011101000",
						 "001010000001110100010000",
						 "001010000001110100111000",
						 "001010000001110101100000",
						 "001010000001101100001000",
						 "001010000001101100110000",
						 "001010000001101101011000",
						 "001010000001101110000000",
						 "001010000001101110101000",
						 "001010000001101111010000",
						 "001010000001101111111000",
						 "001010000001110000100000",
						 "001010000001110001001000",
						 "001010000001110001110000",
						 "001010000001110010011000",
						 "001010000001110011000000",
						 "001010000001110011101000",
						 "001010000001110100010000",
						 "001010000001110100111000",
						 "001010000001110101100000",
						 "001010000001101100001000",
						 "001010000001101100101111",
						 "001010000001101101010110",
						 "001010000001101101111101",
						 "001010000001101110100100",
						 "001010000001101111001011",
						 "001010000001101111110010",
						 "001010000001110000011001",
						 "001010000001110001000000",
						 "001010000001110001100111",
						 "001010000001110010001110",
						 "001010000001110010110101",
						 "001010000001110011011100",
						 "001010000001110100000011",
						 "001010000001110100101010",
						 "001010000001110101010001",
						 "001010000001101100001000",
						 "001010000001101100101111",
						 "001010000001101101010110",
						 "001010000001101101111101",
						 "001010000001101110100100",
						 "001010000001101111001011",
						 "001010000001101111110010",
						 "001010000001110000011001",
						 "001010000001110001000000",
						 "001010000001110001100111",
						 "001010000001110010001110",
						 "001010000001110010110101",
						 "001010000001110011011100",
						 "001010000001110100000011",
						 "001010000001110100101010",
						 "001010000001110101010001",
						 "001010000001101100001000",
						 "001010000001101100101110",
						 "001010000001101101010100",
						 "001010000001101101111010",
						 "001010000001101110100000",
						 "001010000001101111000110",
						 "001010000001101111101100",
						 "001010000001110000010010",
						 "001010000001110000111000",
						 "001010000001110001011110",
						 "001010000001110010000100",
						 "001010000001110010101010",
						 "001010000001110011010000",
						 "001010000001110011110110",
						 "001010000001110100011100",
						 "001010000001110101000010",
						 "001010000001101100001000",
						 "001010000001101100101110",
						 "001010000001101101010100",
						 "001010000001101101111010",
						 "001010000001101110100000",
						 "001010000001101111000110",
						 "001010000001101111101100",
						 "001010000001110000010010",
						 "001010000001110000111000",
						 "001010000001110001011110",
						 "001010000001110010000100",
						 "001010000001110010101010",
						 "001010000001110011010000",
						 "001010000001110011110110",
						 "001010000001110100011100",
						 "001010000001110101000010",
						 "001010000001101100001000",
						 "001010000001101100101110",
						 "001010000001101101010100",
						 "001010000001101101111010",
						 "001010000001101110100000",
						 "001010000001101111000110",
						 "001010000001101111101100",
						 "001010000001110000010010",
						 "001010000001110000111000",
						 "001010000001110001011110",
						 "001010000001110010000100",
						 "001010000001110010101010",
						 "001010000001110011010000",
						 "001010000001110011110110",
						 "001010000001110100011100",
						 "001010000001110101000010",
						 "001010000001101100001000",
						 "001010000001101100101101",
						 "001010000001101101010010",
						 "001010000001101101110111",
						 "001010000001101110011100",
						 "001010000001101111000001",
						 "001010000001101111100110",
						 "001010000001110000001011",
						 "001010000001110000110000",
						 "001010000001110001010101",
						 "001010000001110001111010",
						 "001010000001110010011111",
						 "001010000001110011000100",
						 "001010000001110011101001",
						 "001010000001110100001110",
						 "001010000001110100110011",
						 "001010000001101100001000",
						 "001010000001101100101101",
						 "001010000001101101010010",
						 "001010000001101101110111",
						 "001010000001101110011100",
						 "001010000001101111000001",
						 "001010000001101111100110",
						 "001010000001110000001011",
						 "001010000001110000110000",
						 "001010000001110001010101",
						 "001010000001110001111010",
						 "001010000001110010011111",
						 "001010000001110011000100",
						 "001010000001110011101001",
						 "001010000001110100001110",
						 "001010000001110100110011",
						 "001010000001101100001000",
						 "001010000001101100101100",
						 "001010000001101101010000",
						 "001010000001101101110100",
						 "001010000001101110011000",
						 "001010000001101110111100",
						 "001010000001101111100000",
						 "001010000001110000000100",
						 "001010000001110000101000",
						 "001010000001110001001100",
						 "001010000001110001110000",
						 "001010000001110010010100",
						 "001010000001110010111000",
						 "001010000001110011011100",
						 "001010000001110100000000",
						 "001010000001110100100100",
						 "001010000001101100001000",
						 "001010000001101100101100",
						 "001010000001101101010000",
						 "001010000001101101110100",
						 "001010000001101110011000",
						 "001010000001101110111100",
						 "001010000001101111100000",
						 "001010000001110000000100",
						 "001010000001110000101000",
						 "001010000001110001001100",
						 "001010000001110001110000",
						 "001010000001110010010100",
						 "001010000001110010111000",
						 "001010000001110011011100",
						 "001010000001110100000000",
						 "001010000001110100100100",
						 "001010000001101100001000",
						 "001010000001101100101100",
						 "001010000001101101010000",
						 "001010000001101101110100",
						 "001010000001101110011000",
						 "001010000001101110111100",
						 "001010000001101111100000",
						 "001010000001110000000100",
						 "001010000001110000101000",
						 "001010000001110001001100",
						 "001010000001110001110000",
						 "001010000001110010010100",
						 "001010000001110010111000",
						 "001010000001110011011100",
						 "001010000001110100000000",
						 "001010000001110100100100",
						 "001010000100001111000110",
						 "001010000100001111101001",
						 "001010000100010000001100",
						 "001010000100010000101111",
						 "001010000100010001010010",
						 "001010000100010001110101",
						 "001010000100010010011000",
						 "001010000100010010111011",
						 "001010000100010011011110",
						 "001010000100010100000001",
						 "001010000100010100100100",
						 "001010000100010101000111",
						 "001010000100010101101010",
						 "001010000100010110001101",
						 "001010000100010110110000",
						 "001010000100010111010011",
						 "001010000100001111000110",
						 "001010000100001111101001",
						 "001010000100010000001100",
						 "001010000100010000101111",
						 "001010000100010001010010",
						 "001010000100010001110101",
						 "001010000100010010011000",
						 "001010000100010010111011",
						 "001010000100010011011110",
						 "001010000100010100000001",
						 "001010000100010100100100",
						 "001010000100010101000111",
						 "001010000100010101101010",
						 "001010000100010110001101",
						 "001010000100010110110000",
						 "001010000100010111010011",
						 "001010000100001111000110",
						 "001010000100001111101001",
						 "001010000100010000001100",
						 "001010000100010000101111",
						 "001010000100010001010010",
						 "001010000100010001110101",
						 "001010000100010010011000",
						 "001010000100010010111011",
						 "001010000100010011011110",
						 "001010000100010100000001",
						 "001010000100010100100100",
						 "001010000100010101000111",
						 "001010000100010101101010",
						 "001010000100010110001101",
						 "001010000100010110110000",
						 "001010000100010111010011",
						 "001010000100001111000110",
						 "001010000100001111101000",
						 "001010000100010000001010",
						 "001010000100010000101100",
						 "001010000100010001001110",
						 "001010000100010001110000",
						 "001010000100010010010010",
						 "001010000100010010110100",
						 "001010000100010011010110",
						 "001010000100010011111000",
						 "001010000100010100011010",
						 "001010000100010100111100",
						 "001010000100010101011110",
						 "001010000100010110000000",
						 "001010000100010110100010",
						 "001010000100010111000100",
						 "001010000100001111000110",
						 "001010000100001111101000",
						 "001010000100010000001010",
						 "001010000100010000101100",
						 "001010000100010001001110",
						 "001010000100010001110000",
						 "001010000100010010010010",
						 "001010000100010010110100",
						 "001010000100010011010110",
						 "001010000100010011111000",
						 "001010000100010100011010",
						 "001010000100010100111100",
						 "001010000100010101011110",
						 "001010000100010110000000",
						 "001010000100010110100010",
						 "001010000100010111000100",
						 "001010000100001111000110",
						 "001010000100001111100111",
						 "001010000100010000001000",
						 "001010000100010000101001",
						 "001010000100010001001010",
						 "001010000100010001101011",
						 "001010000100010010001100",
						 "001010000100010010101101",
						 "001010000100010011001110",
						 "001010000100010011101111",
						 "001010000100010100010000",
						 "001010000100010100110001",
						 "001010000100010101010010",
						 "001010000100010101110011",
						 "001010000100010110010100",
						 "001010000100010110110101",
						 "001010000100001111000110",
						 "001010000100001111100111",
						 "001010000100010000001000",
						 "001010000100010000101001",
						 "001010000100010001001010",
						 "001010000100010001101011",
						 "001010000100010010001100",
						 "001010000100010010101101",
						 "001010000100010011001110",
						 "001010000100010011101111",
						 "001010000100010100010000",
						 "001010000100010100110001",
						 "001010000100010101010010",
						 "001010000100010101110011",
						 "001010000100010110010100",
						 "001010000100010110110101",
						 "001010000100001111000110",
						 "001010000100001111100111",
						 "001010000100010000001000",
						 "001010000100010000101001",
						 "001010000100010001001010",
						 "001010000100010001101011",
						 "001010000100010010001100",
						 "001010000100010010101101",
						 "001010000100010011001110",
						 "001010000100010011101111",
						 "001010000100010100010000",
						 "001010000100010100110001",
						 "001010000100010101010010",
						 "001010000100010101110011",
						 "001010000100010110010100",
						 "001010000100010110110101",
						 "001010000100001111000110",
						 "001010000100001111100110",
						 "001010000100010000000110",
						 "001010000100010000100110",
						 "001010000100010001000110",
						 "001010000100010001100110",
						 "001010000100010010000110",
						 "001010000100010010100110",
						 "001010000100010011000110",
						 "001010000100010011100110",
						 "001010000100010100000110",
						 "001010000100010100100110",
						 "001010000100010101000110",
						 "001010000100010101100110",
						 "001010000100010110000110",
						 "001010000100010110100110",
						 "001010000100001111000110",
						 "001010000100001111100110",
						 "001010000100010000000110",
						 "001010000100010000100110",
						 "001010000100010001000110",
						 "001010000100010001100110",
						 "001010000100010010000110",
						 "001010000100010010100110",
						 "001010000100010011000110",
						 "001010000100010011100110",
						 "001010000100010100000110",
						 "001010000100010100100110",
						 "001010000100010101000110",
						 "001010000100010101100110",
						 "001010000100010110000110",
						 "001010000100010110100110",
						 "001010000100001111000110",
						 "001010000100001111100101",
						 "001010000100010000000100",
						 "001010000100010000100011",
						 "001010000100010001000010",
						 "001010000100010001100001",
						 "001010000100010010000000",
						 "001010000100010010011111",
						 "001010000100010010111110",
						 "001010000100010011011101",
						 "001010000100010011111100",
						 "001010000100010100011011",
						 "001010000100010100111010",
						 "001010000100010101011001",
						 "001010000100010101111000",
						 "001010000100010110010111",
						 "001010000100001111000110",
						 "001010000100001111100101",
						 "001010000100010000000100",
						 "001010000100010000100011",
						 "001010000100010001000010",
						 "001010000100010001100001",
						 "001010000100010010000000",
						 "001010000100010010011111",
						 "001010000100010010111110",
						 "001010000100010011011101",
						 "001010000100010011111100",
						 "001010000100010100011011",
						 "001010000100010100111010",
						 "001010000100010101011001",
						 "001010000100010101111000",
						 "001010000100010110010111",
						 "001010000100001111000110",
						 "001010000100001111100101",
						 "001010000100010000000100",
						 "001010000100010000100011",
						 "001010000100010001000010",
						 "001010000100010001100001",
						 "001010000100010010000000",
						 "001010000100010010011111",
						 "001010000100010010111110",
						 "001010000100010011011101",
						 "001010000100010011111100",
						 "001010000100010100011011",
						 "001010000100010100111010",
						 "001010000100010101011001",
						 "001010000100010101111000",
						 "001010000100010110010111",
						 "001010000100001111000110",
						 "001010000100001111100100",
						 "001010000100010000000010",
						 "001010000100010000100000",
						 "001010000100010000111110",
						 "001010000100010001011100",
						 "001010000100010001111010",
						 "001010000100010010011000",
						 "001010000100010010110110",
						 "001010000100010011010100",
						 "001010000100010011110010",
						 "001010000100010100010000",
						 "001010000100010100101110",
						 "001010000100010101001100",
						 "001010000100010101101010",
						 "001010000100010110001000",
						 "001010000100001111000110",
						 "001010000100001111100100",
						 "001010000100010000000010",
						 "001010000100010000100000",
						 "001010000100010000111110",
						 "001010000100010001011100",
						 "001010000100010001111010",
						 "001010000100010010011000",
						 "001010000100010010110110",
						 "001010000100010011010100",
						 "001010000100010011110010",
						 "001010000100010100010000",
						 "001010000100010100101110",
						 "001010000100010101001100",
						 "001010000100010101101010",
						 "001010000100010110001000",
						 "001010000100001111000110",
						 "001010000100001111100011",
						 "001010000100010000000000",
						 "001010000100010000011101",
						 "001010000100010000111010",
						 "001010000100010001010111",
						 "001010000100010001110100",
						 "001010000100010010010001",
						 "001010000100010010101110",
						 "001010000100010011001011",
						 "001010000100010011101000",
						 "001010000100010100000101",
						 "001010000100010100100010",
						 "001010000100010100111111",
						 "001010000100010101011100",
						 "001010000100010101111001",
						 "001010000100001111000110",
						 "001010000100001111100011",
						 "001010000100010000000000",
						 "001010000100010000011101",
						 "001010000100010000111010",
						 "001010000100010001010111",
						 "001010000100010001110100",
						 "001010000100010010010001",
						 "001010000100010010101110",
						 "001010000100010011001011",
						 "001010000100010011101000",
						 "001010000100010100000101",
						 "001010000100010100100010",
						 "001010000100010100111111",
						 "001010000100010101011100",
						 "001010000100010101111001",
						 "001010000100001111000110",
						 "001010000100001111100011",
						 "001010000100010000000000",
						 "001010000100010000011101",
						 "001010000100010000111010",
						 "001010000100010001010111",
						 "001010000100010001110100",
						 "001010000100010010010001",
						 "001010000100010010101110",
						 "001010000100010011001011",
						 "001010000100010011101000",
						 "001010000100010100000101",
						 "001010000100010100100010",
						 "001010000100010100111111",
						 "001010000100010101011100",
						 "001010000100010101111001",
						 "001010000100001111000110",
						 "001010000100001111100010",
						 "001010000100001111111110",
						 "001010000100010000011010",
						 "001010000100010000110110",
						 "001010000100010001010010",
						 "001010000100010001101110",
						 "001010000100010010001010",
						 "001010000100010010100110",
						 "001010000100010011000010",
						 "001010000100010011011110",
						 "001010000100010011111010",
						 "001010000100010100010110",
						 "001010000100010100110010",
						 "001010000100010101001110",
						 "001010000100010101101010",
						 "001010000100001111000110",
						 "001010000100001111100010",
						 "001010000100001111111110",
						 "001010000100010000011010",
						 "001010000100010000110110",
						 "001010000100010001010010",
						 "001010000100010001101110",
						 "001010000100010010001010",
						 "001010000100010010100110",
						 "001010000100010011000010",
						 "001010000100010011011110",
						 "001010000100010011111010",
						 "001010000100010100010110",
						 "001010000100010100110010",
						 "001010000100010101001110",
						 "001010000100010101101010",
						 "001010000100001111000110",
						 "001010000100001111100010",
						 "001010000100001111111110",
						 "001010000100010000011010",
						 "001010000100010000110110",
						 "001010000100010001010010",
						 "001010000100010001101110",
						 "001010000100010010001010",
						 "001010000100010010100110",
						 "001010000100010011000010",
						 "001010000100010011011110",
						 "001010000100010011111010",
						 "001010000100010100010110",
						 "001010000100010100110010",
						 "001010000100010101001110",
						 "001010000100010101101010",
						 "001010000110110010000100",
						 "001010000110110010011111",
						 "001010000110110010111010",
						 "001010000110110011010101",
						 "001010000110110011110000",
						 "001010000110110100001011",
						 "001010000110110100100110",
						 "001010000110110101000001",
						 "001010000110110101011100",
						 "001010000110110101110111",
						 "001010000110110110010010",
						 "001010000110110110101101",
						 "001010000110110111001000",
						 "001010000110110111100011",
						 "001010000110110111111110",
						 "001010000110111000011001",
						 "001010000110110010000100",
						 "001010000110110010011111",
						 "001010000110110010111010",
						 "001010000110110011010101",
						 "001010000110110011110000",
						 "001010000110110100001011",
						 "001010000110110100100110",
						 "001010000110110101000001",
						 "001010000110110101011100",
						 "001010000110110101110111",
						 "001010000110110110010010",
						 "001010000110110110101101",
						 "001010000110110111001000",
						 "001010000110110111100011",
						 "001010000110110111111110",
						 "001010000110111000011001",
						 "001010000110110010000100",
						 "001010000110110010011110",
						 "001010000110110010111000",
						 "001010000110110011010010",
						 "001010000110110011101100",
						 "001010000110110100000110",
						 "001010000110110100100000",
						 "001010000110110100111010",
						 "001010000110110101010100",
						 "001010000110110101101110",
						 "001010000110110110001000",
						 "001010000110110110100010",
						 "001010000110110110111100",
						 "001010000110110111010110",
						 "001010000110110111110000",
						 "001010000110111000001010",
						 "001010000110110010000100",
						 "001010000110110010011110",
						 "001010000110110010111000",
						 "001010000110110011010010",
						 "001010000110110011101100",
						 "001010000110110100000110",
						 "001010000110110100100000",
						 "001010000110110100111010",
						 "001010000110110101010100",
						 "001010000110110101101110",
						 "001010000110110110001000",
						 "001010000110110110100010",
						 "001010000110110110111100",
						 "001010000110110111010110",
						 "001010000110110111110000",
						 "001010000110111000001010",
						 "001010000110110010000100",
						 "001010000110110010011110",
						 "001010000110110010111000",
						 "001010000110110011010010",
						 "001010000110110011101100",
						 "001010000110110100000110",
						 "001010000110110100100000",
						 "001010000110110100111010",
						 "001010000110110101010100",
						 "001010000110110101101110",
						 "001010000110110110001000",
						 "001010000110110110100010",
						 "001010000110110110111100",
						 "001010000110110111010110",
						 "001010000110110111110000",
						 "001010000110111000001010",
						 "001010000110110010000100",
						 "001010000110110010011101",
						 "001010000110110010110110",
						 "001010000110110011001111",
						 "001010000110110011101000",
						 "001010000110110100000001",
						 "001010000110110100011010",
						 "001010000110110100110011",
						 "001010000110110101001100",
						 "001010000110110101100101",
						 "001010000110110101111110",
						 "001010000110110110010111",
						 "001010000110110110110000",
						 "001010000110110111001001",
						 "001010000110110111100010",
						 "001010000110110111111011",
						 "001010000110110010000100",
						 "001010000110110010011101",
						 "001010000110110010110110",
						 "001010000110110011001111",
						 "001010000110110011101000",
						 "001010000110110100000001",
						 "001010000110110100011010",
						 "001010000110110100110011",
						 "001010000110110101001100",
						 "001010000110110101100101",
						 "001010000110110101111110",
						 "001010000110110110010111",
						 "001010000110110110110000",
						 "001010000110110111001001",
						 "001010000110110111100010",
						 "001010000110110111111011",
						 "001010000110110010000100",
						 "001010000110110010011100",
						 "001010000110110010110100",
						 "001010000110110011001100",
						 "001010000110110011100100",
						 "001010000110110011111100",
						 "001010000110110100010100",
						 "001010000110110100101100",
						 "001010000110110101000100",
						 "001010000110110101011100",
						 "001010000110110101110100",
						 "001010000110110110001100",
						 "001010000110110110100100",
						 "001010000110110110111100",
						 "001010000110110111010100",
						 "001010000110110111101100",
						 "001010000110110010000100",
						 "001010000110110010011100",
						 "001010000110110010110100",
						 "001010000110110011001100",
						 "001010000110110011100100",
						 "001010000110110011111100",
						 "001010000110110100010100",
						 "001010000110110100101100",
						 "001010000110110101000100",
						 "001010000110110101011100",
						 "001010000110110101110100",
						 "001010000110110110001100",
						 "001010000110110110100100",
						 "001010000110110110111100",
						 "001010000110110111010100",
						 "001010000110110111101100",
						 "001010000110110010000100",
						 "001010000110110010011100",
						 "001010000110110010110100",
						 "001010000110110011001100",
						 "001010000110110011100100",
						 "001010000110110011111100",
						 "001010000110110100010100",
						 "001010000110110100101100",
						 "001010000110110101000100",
						 "001010000110110101011100",
						 "001010000110110101110100",
						 "001010000110110110001100",
						 "001010000110110110100100",
						 "001010000110110110111100",
						 "001010000110110111010100",
						 "001010000110110111101100",
						 "001010000110110010000100",
						 "001010000110110010011011",
						 "001010000110110010110010",
						 "001010000110110011001001",
						 "001010000110110011100000",
						 "001010000110110011110111",
						 "001010000110110100001110",
						 "001010000110110100100101",
						 "001010000110110100111100",
						 "001010000110110101010011",
						 "001010000110110101101010",
						 "001010000110110110000001",
						 "001010000110110110011000",
						 "001010000110110110101111",
						 "001010000110110111000110",
						 "001010000110110111011101",
						 "001010000110110010000100",
						 "001010000110110010011011",
						 "001010000110110010110010",
						 "001010000110110011001001",
						 "001010000110110011100000",
						 "001010000110110011110111",
						 "001010000110110100001110",
						 "001010000110110100100101",
						 "001010000110110100111100",
						 "001010000110110101010011",
						 "001010000110110101101010",
						 "001010000110110110000001",
						 "001010000110110110011000",
						 "001010000110110110101111",
						 "001010000110110111000110",
						 "001010000110110111011101",
						 "001010000110110010000100",
						 "001010000110110010011010",
						 "001010000110110010110000",
						 "001010000110110011000110",
						 "001010000110110011011100",
						 "001010000110110011110010",
						 "001010000110110100001000",
						 "001010000110110100011110",
						 "001010000110110100110100",
						 "001010000110110101001010",
						 "001010000110110101100000",
						 "001010000110110101110110",
						 "001010000110110110001100",
						 "001010000110110110100010",
						 "001010000110110110111000",
						 "001010000110110111001110",
						 "001010000110110010000100",
						 "001010000110110010011010",
						 "001010000110110010110000",
						 "001010000110110011000110",
						 "001010000110110011011100",
						 "001010000110110011110010",
						 "001010000110110100001000",
						 "001010000110110100011110",
						 "001010000110110100110100",
						 "001010000110110101001010",
						 "001010000110110101100000",
						 "001010000110110101110110",
						 "001010000110110110001100",
						 "001010000110110110100010",
						 "001010000110110110111000",
						 "001010000110110111001110",
						 "001010000110110010000100",
						 "001010000110110010011010",
						 "001010000110110010110000",
						 "001010000110110011000110",
						 "001010000110110011011100",
						 "001010000110110011110010",
						 "001010000110110100001000",
						 "001010000110110100011110",
						 "001010000110110100110100",
						 "001010000110110101001010",
						 "001010000110110101100000",
						 "001010000110110101110110",
						 "001010000110110110001100",
						 "001010000110110110100010",
						 "001010000110110110111000",
						 "001010000110110111001110",
						 "001010000110110010000100",
						 "001010000110110010011001",
						 "001010000110110010101110",
						 "001010000110110011000011",
						 "001010000110110011011000",
						 "001010000110110011101101",
						 "001010000110110100000010",
						 "001010000110110100010111",
						 "001010000110110100101100",
						 "001010000110110101000001",
						 "001010000110110101010110",
						 "001010000110110101101011",
						 "001010000110110110000000",
						 "001010000110110110010101",
						 "001010000110110110101010",
						 "001010000110110110111111",
						 "001010000110110010000100",
						 "001010000110110010011001",
						 "001010000110110010101110",
						 "001010000110110011000011",
						 "001010000110110011011000",
						 "001010000110110011101101",
						 "001010000110110100000010",
						 "001010000110110100010111",
						 "001010000110110100101100",
						 "001010000110110101000001",
						 "001010000110110101010110",
						 "001010000110110101101011",
						 "001010000110110110000000",
						 "001010000110110110010101",
						 "001010000110110110101010",
						 "001010000110110110111111",
						 "001010000110110010000100",
						 "001010000110110010011001",
						 "001010000110110010101110",
						 "001010000110110011000011",
						 "001010000110110011011000",
						 "001010000110110011101101",
						 "001010000110110100000010",
						 "001010000110110100010111",
						 "001010000110110100101100",
						 "001010000110110101000001",
						 "001010000110110101010110",
						 "001010000110110101101011",
						 "001010000110110110000000",
						 "001010000110110110010101",
						 "001010000110110110101010",
						 "001010000110110110111111",
						 "001010000110110010000100",
						 "001010000110110010011000",
						 "001010000110110010101100",
						 "001010000110110011000000",
						 "001010000110110011010100",
						 "001010000110110011101000",
						 "001010000110110011111100",
						 "001010000110110100010000",
						 "001010000110110100100100",
						 "001010000110110100111000",
						 "001010000110110101001100",
						 "001010000110110101100000",
						 "001010000110110101110100",
						 "001010000110110110001000",
						 "001010000110110110011100",
						 "001010000110110110110000",
						 "001010000110110010000100",
						 "001010000110110010011000",
						 "001010000110110010101100",
						 "001010000110110011000000",
						 "001010000110110011010100",
						 "001010000110110011101000",
						 "001010000110110011111100",
						 "001010000110110100010000",
						 "001010000110110100100100",
						 "001010000110110100111000",
						 "001010000110110101001100",
						 "001010000110110101100000",
						 "001010000110110101110100",
						 "001010000110110110001000",
						 "001010000110110110011100",
						 "001010000110110110110000",
						 "001010000110110010000100",
						 "001010000110110010010111",
						 "001010000110110010101010",
						 "001010000110110010111101",
						 "001010000110110011010000",
						 "001010000110110011100011",
						 "001010000110110011110110",
						 "001010000110110100001001",
						 "001010000110110100011100",
						 "001010000110110100101111",
						 "001010000110110101000010",
						 "001010000110110101010101",
						 "001010000110110101101000",
						 "001010000110110101111011",
						 "001010000110110110001110",
						 "001010000110110110100001",
						 "001010000110110010000100",
						 "001010000110110010010111",
						 "001010000110110010101010",
						 "001010000110110010111101",
						 "001010000110110011010000",
						 "001010000110110011100011",
						 "001010000110110011110110",
						 "001010000110110100001001",
						 "001010000110110100011100",
						 "001010000110110100101111",
						 "001010000110110101000010",
						 "001010000110110101010101",
						 "001010000110110101101000",
						 "001010000110110101111011",
						 "001010000110110110001110",
						 "001010000110110110100001",
						 "001010000110110010000100",
						 "001010000110110010010111",
						 "001010000110110010101010",
						 "001010000110110010111101",
						 "001010000110110011010000",
						 "001010000110110011100011",
						 "001010000110110011110110",
						 "001010000110110100001001",
						 "001010000110110100011100",
						 "001010000110110100101111",
						 "001010000110110101000010",
						 "001010000110110101010101",
						 "001010000110110101101000",
						 "001010000110110101111011",
						 "001010000110110110001110",
						 "001010000110110110100001",
						 "001010000110110010000100",
						 "001010000110110010010110",
						 "001010000110110010101000",
						 "001010000110110010111010",
						 "001010000110110011001100",
						 "001010000110110011011110",
						 "001010000110110011110000",
						 "001010000110110100000010",
						 "001010000110110100010100",
						 "001010000110110100100110",
						 "001010000110110100111000",
						 "001010000110110101001010",
						 "001010000110110101011100",
						 "001010000110110101101110",
						 "001010000110110110000000",
						 "001010000110110110010010",
						 "001010000110110010000100",
						 "001010000110110010010110",
						 "001010000110110010101000",
						 "001010000110110010111010",
						 "001010000110110011001100",
						 "001010000110110011011110",
						 "001010000110110011110000",
						 "001010000110110100000010",
						 "001010000110110100010100",
						 "001010000110110100100110",
						 "001010000110110100111000",
						 "001010000110110101001010",
						 "001010000110110101011100",
						 "001010000110110101101110",
						 "001010000110110110000000",
						 "001010000110110110010010",
						 "001010000110110010000100",
						 "001010000110110010010101",
						 "001010000110110010100110",
						 "001010000110110010110111",
						 "001010000110110011001000",
						 "001010000110110011011001",
						 "001010000110110011101010",
						 "001010000110110011111011",
						 "001010000110110100001100",
						 "001010000110110100011101",
						 "001010000110110100101110",
						 "001010000110110100111111",
						 "001010000110110101010000",
						 "001010000110110101100001",
						 "001010000110110101110010",
						 "001010000110110110000011",
						 "001010000110110010000100",
						 "001010000110110010010101",
						 "001010000110110010100110",
						 "001010000110110010110111",
						 "001010000110110011001000",
						 "001010000110110011011001",
						 "001010000110110011101010",
						 "001010000110110011111011",
						 "001010000110110100001100",
						 "001010000110110100011101",
						 "001010000110110100101110",
						 "001010000110110100111111",
						 "001010000110110101010000",
						 "001010000110110101100001",
						 "001010000110110101110010",
						 "001010000110110110000011",
						 "001010000110110010000100",
						 "001010000110110010010101",
						 "001010000110110010100110",
						 "001010000110110010110111",
						 "001010000110110011001000",
						 "001010000110110011011001",
						 "001010000110110011101010",
						 "001010000110110011111011",
						 "001010000110110100001100",
						 "001010000110110100011101",
						 "001010000110110100101110",
						 "001010000110110100111111",
						 "001010000110110101010000",
						 "001010000110110101100001",
						 "001010000110110101110010",
						 "001010000110110110000011",
						 "001010000110110010000100",
						 "001010000110110010010100",
						 "001010000110110010100100",
						 "001010000110110010110100",
						 "001010000110110011000100",
						 "001010000110110011010100",
						 "001010000110110011100100",
						 "001010000110110011110100",
						 "001010000110110100000100",
						 "001010000110110100010100",
						 "001010000110110100100100",
						 "001010000110110100110100",
						 "001010000110110101000100",
						 "001010000110110101010100",
						 "001010000110110101100100",
						 "001010000110110101110100",
						 "001010000110110010000100",
						 "001010000110110010010100",
						 "001010000110110010100100",
						 "001010000110110010110100",
						 "001010000110110011000100",
						 "001010000110110011010100",
						 "001010000110110011100100",
						 "001010000110110011110100",
						 "001010000110110100000100",
						 "001010000110110100010100",
						 "001010000110110100100100",
						 "001010000110110100110100",
						 "001010000110110101000100",
						 "001010000110110101010100",
						 "001010000110110101100100",
						 "001010000110110101110100",
						 "001010001001010101000010",
						 "001010001001010101010001",
						 "001010001001010101100000",
						 "001010001001010101101111",
						 "001010001001010101111110",
						 "001010001001010110001101",
						 "001010001001010110011100",
						 "001010001001010110101011",
						 "001010001001010110111010",
						 "001010001001010111001001",
						 "001010001001010111011000",
						 "001010001001010111100111",
						 "001010001001010111110110",
						 "001010001001011000000101",
						 "001010001001011000010100",
						 "001010001001011000100011",
						 "001010001001010101000010",
						 "001010001001010101010001",
						 "001010001001010101100000",
						 "001010001001010101101111",
						 "001010001001010101111110",
						 "001010001001010110001101",
						 "001010001001010110011100",
						 "001010001001010110101011",
						 "001010001001010110111010",
						 "001010001001010111001001",
						 "001010001001010111011000",
						 "001010001001010111100111",
						 "001010001001010111110110",
						 "001010001001011000000101",
						 "001010001001011000010100",
						 "001010001001011000100011",
						 "001010001001010101000010",
						 "001010001001010101010001",
						 "001010001001010101100000",
						 "001010001001010101101111",
						 "001010001001010101111110",
						 "001010001001010110001101",
						 "001010001001010110011100",
						 "001010001001010110101011",
						 "001010001001010110111010",
						 "001010001001010111001001",
						 "001010001001010111011000",
						 "001010001001010111100111",
						 "001010001001010111110110",
						 "001010001001011000000101",
						 "001010001001011000010100",
						 "001010001001011000100011",
						 "001010001001010101000010",
						 "001010001001010101010000",
						 "001010001001010101011110",
						 "001010001001010101101100",
						 "001010001001010101111010",
						 "001010001001010110001000",
						 "001010001001010110010110",
						 "001010001001010110100100",
						 "001010001001010110110010",
						 "001010001001010111000000",
						 "001010001001010111001110",
						 "001010001001010111011100",
						 "001010001001010111101010",
						 "001010001001010111111000",
						 "001010001001011000000110",
						 "001010001001011000010100",
						 "001010001001010101000010",
						 "001010001001010101010000",
						 "001010001001010101011110",
						 "001010001001010101101100",
						 "001010001001010101111010",
						 "001010001001010110001000",
						 "001010001001010110010110",
						 "001010001001010110100100",
						 "001010001001010110110010",
						 "001010001001010111000000",
						 "001010001001010111001110",
						 "001010001001010111011100",
						 "001010001001010111101010",
						 "001010001001010111111000",
						 "001010001001011000000110",
						 "001010001001011000010100",
						 "001010001001010101000010",
						 "001010001001010101001111",
						 "001010001001010101011100",
						 "001010001001010101101001",
						 "001010001001010101110110",
						 "001010001001010110000011",
						 "001010001001010110010000",
						 "001010001001010110011101",
						 "001010001001010110101010",
						 "001010001001010110110111",
						 "001010001001010111000100",
						 "001010001001010111010001",
						 "001010001001010111011110",
						 "001010001001010111101011",
						 "001010001001010111111000",
						 "001010001001011000000101",
						 "001010001001010101000010",
						 "001010001001010101001111",
						 "001010001001010101011100",
						 "001010001001010101101001",
						 "001010001001010101110110",
						 "001010001001010110000011",
						 "001010001001010110010000",
						 "001010001001010110011101",
						 "001010001001010110101010",
						 "001010001001010110110111",
						 "001010001001010111000100",
						 "001010001001010111010001",
						 "001010001001010111011110",
						 "001010001001010111101011",
						 "001010001001010111111000",
						 "001010001001011000000101",
						 "001010001001010101000010",
						 "001010001001010101001111",
						 "001010001001010101011100",
						 "001010001001010101101001",
						 "001010001001010101110110",
						 "001010001001010110000011",
						 "001010001001010110010000",
						 "001010001001010110011101",
						 "001010001001010110101010",
						 "001010001001010110110111",
						 "001010001001010111000100",
						 "001010001001010111010001",
						 "001010001001010111011110",
						 "001010001001010111101011",
						 "001010001001010111111000",
						 "001010001001011000000101",
						 "001010001001010101000010",
						 "001010001001010101001110",
						 "001010001001010101011010",
						 "001010001001010101100110",
						 "001010001001010101110010",
						 "001010001001010101111110",
						 "001010001001010110001010",
						 "001010001001010110010110",
						 "001010001001010110100010",
						 "001010001001010110101110",
						 "001010001001010110111010",
						 "001010001001010111000110",
						 "001010001001010111010010",
						 "001010001001010111011110",
						 "001010001001010111101010",
						 "001010001001010111110110",
						 "001010001001010101000010",
						 "001010001001010101001110",
						 "001010001001010101011010",
						 "001010001001010101100110",
						 "001010001001010101110010",
						 "001010001001010101111110",
						 "001010001001010110001010",
						 "001010001001010110010110",
						 "001010001001010110100010",
						 "001010001001010110101110",
						 "001010001001010110111010",
						 "001010001001010111000110",
						 "001010001001010111010010",
						 "001010001001010111011110",
						 "001010001001010111101010",
						 "001010001001010111110110",
						 "001010001001010101000010",
						 "001010001001010101001110",
						 "001010001001010101011010",
						 "001010001001010101100110",
						 "001010001001010101110010",
						 "001010001001010101111110",
						 "001010001001010110001010",
						 "001010001001010110010110",
						 "001010001001010110100010",
						 "001010001001010110101110",
						 "001010001001010110111010",
						 "001010001001010111000110",
						 "001010001001010111010010",
						 "001010001001010111011110",
						 "001010001001010111101010",
						 "001010001001010111110110",
						 "001010001001010101000010",
						 "001010001001010101001101",
						 "001010001001010101011000",
						 "001010001001010101100011",
						 "001010001001010101101110",
						 "001010001001010101111001",
						 "001010001001010110000100",
						 "001010001001010110001111",
						 "001010001001010110011010",
						 "001010001001010110100101",
						 "001010001001010110110000",
						 "001010001001010110111011",
						 "001010001001010111000110",
						 "001010001001010111010001",
						 "001010001001010111011100",
						 "001010001001010111100111",
						 "001010001001010101000010",
						 "001010001001010101001101",
						 "001010001001010101011000",
						 "001010001001010101100011",
						 "001010001001010101101110",
						 "001010001001010101111001",
						 "001010001001010110000100",
						 "001010001001010110001111",
						 "001010001001010110011010",
						 "001010001001010110100101",
						 "001010001001010110110000",
						 "001010001001010110111011",
						 "001010001001010111000110",
						 "001010001001010111010001",
						 "001010001001010111011100",
						 "001010001001010111100111",
						 "001010001001010101000010",
						 "001010001001010101001100",
						 "001010001001010101010110",
						 "001010001001010101100000",
						 "001010001001010101101010",
						 "001010001001010101110100",
						 "001010001001010101111110",
						 "001010001001010110001000",
						 "001010001001010110010010",
						 "001010001001010110011100",
						 "001010001001010110100110",
						 "001010001001010110110000",
						 "001010001001010110111010",
						 "001010001001010111000100",
						 "001010001001010111001110",
						 "001010001001010111011000",
						 "001010001001010101000010",
						 "001010001001010101001100",
						 "001010001001010101010110",
						 "001010001001010101100000",
						 "001010001001010101101010",
						 "001010001001010101110100",
						 "001010001001010101111110",
						 "001010001001010110001000",
						 "001010001001010110010010",
						 "001010001001010110011100",
						 "001010001001010110100110",
						 "001010001001010110110000",
						 "001010001001010110111010",
						 "001010001001010111000100",
						 "001010001001010111001110",
						 "001010001001010111011000",
						 "001010001001010101000010",
						 "001010001001010101001100",
						 "001010001001010101010110",
						 "001010001001010101100000",
						 "001010001001010101101010",
						 "001010001001010101110100",
						 "001010001001010101111110",
						 "001010001001010110001000",
						 "001010001001010110010010",
						 "001010001001010110011100",
						 "001010001001010110100110",
						 "001010001001010110110000",
						 "001010001001010110111010",
						 "001010001001010111000100",
						 "001010001001010111001110",
						 "001010001001010111011000",
						 "001010001001010101000010",
						 "001010001001010101001011",
						 "001010001001010101010100",
						 "001010001001010101011101",
						 "001010001001010101100110",
						 "001010001001010101101111",
						 "001010001001010101111000",
						 "001010001001010110000001",
						 "001010001001010110001010",
						 "001010001001010110010011",
						 "001010001001010110011100",
						 "001010001001010110100101",
						 "001010001001010110101110",
						 "001010001001010110110111",
						 "001010001001010111000000",
						 "001010001001010111001001",
						 "001010001001010101000010",
						 "001010001001010101001011",
						 "001010001001010101010100",
						 "001010001001010101011101",
						 "001010001001010101100110",
						 "001010001001010101101111",
						 "001010001001010101111000",
						 "001010001001010110000001",
						 "001010001001010110001010",
						 "001010001001010110010011",
						 "001010001001010110011100",
						 "001010001001010110100101",
						 "001010001001010110101110",
						 "001010001001010110110111",
						 "001010001001010111000000",
						 "001010001001010111001001",
						 "001010001001010101000010",
						 "001010001001010101001010",
						 "001010001001010101010010",
						 "001010001001010101011010",
						 "001010001001010101100010",
						 "001010001001010101101010",
						 "001010001001010101110010",
						 "001010001001010101111010",
						 "001010001001010110000010",
						 "001010001001010110001010",
						 "001010001001010110010010",
						 "001010001001010110011010",
						 "001010001001010110100010",
						 "001010001001010110101010",
						 "001010001001010110110010",
						 "001010001001010110111010",
						 "001010001001010101000010",
						 "001010001001010101001010",
						 "001010001001010101010010",
						 "001010001001010101011010",
						 "001010001001010101100010",
						 "001010001001010101101010",
						 "001010001001010101110010",
						 "001010001001010101111010",
						 "001010001001010110000010",
						 "001010001001010110001010",
						 "001010001001010110010010",
						 "001010001001010110011010",
						 "001010001001010110100010",
						 "001010001001010110101010",
						 "001010001001010110110010",
						 "001010001001010110111010",
						 "001010001001010101000010",
						 "001010001001010101001010",
						 "001010001001010101010010",
						 "001010001001010101011010",
						 "001010001001010101100010",
						 "001010001001010101101010",
						 "001010001001010101110010",
						 "001010001001010101111010",
						 "001010001001010110000010",
						 "001010001001010110001010",
						 "001010001001010110010010",
						 "001010001001010110011010",
						 "001010001001010110100010",
						 "001010001001010110101010",
						 "001010001001010110110010",
						 "001010001001010110111010",
						 "001010001001010101000010",
						 "001010001001010101001001",
						 "001010001001010101010000",
						 "001010001001010101010111",
						 "001010001001010101011110",
						 "001010001001010101100101",
						 "001010001001010101101100",
						 "001010001001010101110011",
						 "001010001001010101111010",
						 "001010001001010110000001",
						 "001010001001010110001000",
						 "001010001001010110001111",
						 "001010001001010110010110",
						 "001010001001010110011101",
						 "001010001001010110100100",
						 "001010001001010110101011",
						 "001010001001010101000010",
						 "001010001001010101001001",
						 "001010001001010101010000",
						 "001010001001010101010111",
						 "001010001001010101011110",
						 "001010001001010101100101",
						 "001010001001010101101100",
						 "001010001001010101110011",
						 "001010001001010101111010",
						 "001010001001010110000001",
						 "001010001001010110001000",
						 "001010001001010110001111",
						 "001010001001010110010110",
						 "001010001001010110011101",
						 "001010001001010110100100",
						 "001010001001010110101011",
						 "001010001001010101000010",
						 "001010001001010101001000",
						 "001010001001010101001110",
						 "001010001001010101010100",
						 "001010001001010101011010",
						 "001010001001010101100000",
						 "001010001001010101100110",
						 "001010001001010101101100",
						 "001010001001010101110010",
						 "001010001001010101111000",
						 "001010001001010101111110",
						 "001010001001010110000100",
						 "001010001001010110001010",
						 "001010001001010110010000",
						 "001010001001010110010110",
						 "001010001001010110011100",
						 "001010001001010101000010",
						 "001010001001010101001000",
						 "001010001001010101001110",
						 "001010001001010101010100",
						 "001010001001010101011010",
						 "001010001001010101100000",
						 "001010001001010101100110",
						 "001010001001010101101100",
						 "001010001001010101110010",
						 "001010001001010101111000",
						 "001010001001010101111110",
						 "001010001001010110000100",
						 "001010001001010110001010",
						 "001010001001010110010000",
						 "001010001001010110010110",
						 "001010001001010110011100",
						 "001010001001010101000010",
						 "001010001001010101001000",
						 "001010001001010101001110",
						 "001010001001010101010100",
						 "001010001001010101011010",
						 "001010001001010101100000",
						 "001010001001010101100110",
						 "001010001001010101101100",
						 "001010001001010101110010",
						 "001010001001010101111000",
						 "001010001001010101111110",
						 "001010001001010110000100",
						 "001010001001010110001010",
						 "001010001001010110010000",
						 "001010001001010110010110",
						 "001010001001010110011100",
						 "001010001001010101000010",
						 "001010001001010101000111",
						 "001010001001010101001100",
						 "001010001001010101010001",
						 "001010001001010101010110",
						 "001010001001010101011011",
						 "001010001001010101100000",
						 "001010001001010101100101",
						 "001010001001010101101010",
						 "001010001001010101101111",
						 "001010001001010101110100",
						 "001010001001010101111001",
						 "001010001001010101111110",
						 "001010001001010110000011",
						 "001010001001010110001000",
						 "001010001001010110001101",
						 "001010001001010101000010",
						 "001010001001010101000111",
						 "001010001001010101001100",
						 "001010001001010101010001",
						 "001010001001010101010110",
						 "001010001001010101011011",
						 "001010001001010101100000",
						 "001010001001010101100101",
						 "001010001001010101101010",
						 "001010001001010101101111",
						 "001010001001010101110100",
						 "001010001001010101111001",
						 "001010001001010101111110",
						 "001010001001010110000011",
						 "001010001001010110001000",
						 "001010001001010110001101",
						 "001010001001010101000010",
						 "001010001001010101000110",
						 "001010001001010101001010",
						 "001010001001010101001110",
						 "001010001001010101010010",
						 "001010001001010101010110",
						 "001010001001010101011010",
						 "001010001001010101011110",
						 "001010001001010101100010",
						 "001010001001010101100110",
						 "001010001001010101101010",
						 "001010001001010101101110",
						 "001010001001010101110010",
						 "001010001001010101110110",
						 "001010001001010101111010",
						 "001010001001010101111110",
						 "001010001001010101000010",
						 "001010001001010101000110",
						 "001010001001010101001010",
						 "001010001001010101001110",
						 "001010001001010101010010",
						 "001010001001010101010110",
						 "001010001001010101011010",
						 "001010001001010101011110",
						 "001010001001010101100010",
						 "001010001001010101100110",
						 "001010001001010101101010",
						 "001010001001010101101110",
						 "001010001001010101110010",
						 "001010001001010101110110",
						 "001010001001010101111010",
						 "001010001001010101111110",
						 "001010001001010101000010",
						 "001010001001010101000110",
						 "001010001001010101001010",
						 "001010001001010101001110",
						 "001010001001010101010010",
						 "001010001001010101010110",
						 "001010001001010101011010",
						 "001010001001010101011110",
						 "001010001001010101100010",
						 "001010001001010101100110",
						 "001010001001010101101010",
						 "001010001001010101101110",
						 "001010001001010101110010",
						 "001010001001010101110110",
						 "001010001001010101111010",
						 "001010001001010101111110",
						 "001010001001010101000010",
						 "001010001001010101000101",
						 "001010001001010101001000",
						 "001010001001010101001011",
						 "001010001001010101001110",
						 "001010001001010101010001",
						 "001010001001010101010100",
						 "001010001001010101010111",
						 "001010001001010101011010",
						 "001010001001010101011101",
						 "001010001001010101100000",
						 "001010001001010101100011",
						 "001010001001010101100110",
						 "001010001001010101101001",
						 "001010001001010101101100",
						 "001010001001010101101111",
						 "001010001001010101000010",
						 "001010001001010101000101",
						 "001010001001010101001000",
						 "001010001001010101001011",
						 "001010001001010101001110",
						 "001010001001010101010001",
						 "001010001001010101010100",
						 "001010001001010101010111",
						 "001010001001010101011010",
						 "001010001001010101011101",
						 "001010001001010101100000",
						 "001010001001010101100011",
						 "001010001001010101100110",
						 "001010001001010101101001",
						 "001010001001010101101100",
						 "001010001001010101101111",
						 "001010001001010101000010",
						 "001010001001010101000101",
						 "001010001001010101001000",
						 "001010001001010101001011",
						 "001010001001010101001110",
						 "001010001001010101010001",
						 "001010001001010101010100",
						 "001010001001010101010111",
						 "001010001001010101011010",
						 "001010001001010101011101",
						 "001010001001010101100000",
						 "001010001001010101100011",
						 "001010001001010101100110",
						 "001010001001010101101001",
						 "001010001001010101101100",
						 "001010001001010101101111",
						 "001010001001010101000010",
						 "001010001001010101000100",
						 "001010001001010101000110",
						 "001010001001010101001000",
						 "001010001001010101001010",
						 "001010001001010101001100",
						 "001010001001010101001110",
						 "001010001001010101010000",
						 "001010001001010101010010",
						 "001010001001010101010100",
						 "001010001001010101010110",
						 "001010001001010101011000",
						 "001010001001010101011010",
						 "001010001001010101011100",
						 "001010001001010101011110",
						 "001010001001010101100000",
						 "001010001001010101000010",
						 "001010001001010101000100",
						 "001010001001010101000110",
						 "001010001001010101001000",
						 "001010001001010101001010",
						 "001010001001010101001100",
						 "001010001001010101001110",
						 "001010001001010101010000",
						 "001010001001010101010010",
						 "001010001001010101010100",
						 "001010001001010101010110",
						 "001010001001010101011000",
						 "001010001001010101011010",
						 "001010001001010101011100",
						 "001010001001010101011110",
						 "001010001001010101100000",
						 "001010001001010101000010",
						 "001010001001010101000011",
						 "001010001001010101000100",
						 "001010001001010101000101",
						 "001010001001010101000110",
						 "001010001001010101000111",
						 "001010001001010101001000",
						 "001010001001010101001001",
						 "001010001001010101001010",
						 "001010001001010101001011",
						 "001010001001010101001100",
						 "001010001001010101001101",
						 "001010001001010101001110",
						 "001010001001010101001111",
						 "001010001001010101010000",
						 "001010001001010101010001",
						 "001010001001010101000010",
						 "001010001001010101000011",
						 "001010001001010101000100",
						 "001010001001010101000101",
						 "001010001001010101000110",
						 "001010001001010101000111",
						 "001010001001010101001000",
						 "001010001001010101001001",
						 "001010001001010101001010",
						 "001010001001010101001011",
						 "001010001001010101001100",
						 "001010001001010101001101",
						 "001010001001010101001110",
						 "001010001001010101001111",
						 "001010001001010101010000",
						 "001010001001010101010001",
						 "001010001001010101000010",
						 "001010001001010101000011",
						 "001010001001010101000100",
						 "001010001001010101000101",
						 "001010001001010101000110",
						 "001010001001010101000111",
						 "001010001001010101001000",
						 "001010001001010101001001",
						 "001010001001010101001010",
						 "001010001001010101001011",
						 "001010001001010101001100",
						 "001010001001010101001101",
						 "001010001001010101001110",
						 "001010001001010101001111",
						 "001010001001010101010000",
						 "001010001001010101010001",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101000010",
						 "001010001001010101010001",
						 "001010001001010101010000",
						 "001010001001010101001111",
						 "001010001001010101001110",
						 "001010001001010101001101",
						 "001010001001010101001100",
						 "001010001001010101001011",
						 "001010001001010101001010",
						 "001010001001010101001001",
						 "001010001001010101001000",
						 "001010001001010101000111",
						 "001010001001010101000110",
						 "001010001001010101000101",
						 "001010001001010101000100",
						 "001010001001010101000011",
						 "001010001001010101000010",
						 "001010001001010101010001",
						 "001010001001010101010000",
						 "001010001001010101001111",
						 "001010001001010101001110",
						 "001010001001010101001101",
						 "001010001001010101001100",
						 "001010001001010101001011",
						 "001010001001010101001010",
						 "001010001001010101001001",
						 "001010001001010101001000",
						 "001010001001010101000111",
						 "001010001001010101000110",
						 "001010001001010101000101",
						 "001010001001010101000100",
						 "001010001001010101000011",
						 "001010001001010101000010",
						 "001010001001010101010001",
						 "001010001001010101010000",
						 "001010001001010101001111",
						 "001010001001010101001110",
						 "001010001001010101001101",
						 "001010001001010101001100",
						 "001010001001010101001011",
						 "001010001001010101001010",
						 "001010001001010101001001",
						 "001010001001010101001000",
						 "001010001001010101000111",
						 "001010001001010101000110",
						 "001010001001010101000101",
						 "001010001001010101000100",
						 "001010001001010101000011",
						 "001010001001010101000010",
						 "001010001001010101100000",
						 "001010001001010101011110",
						 "001010001001010101011100",
						 "001010001001010101011010",
						 "001010001001010101011000",
						 "001010001001010101010110",
						 "001010001001010101010100",
						 "001010001001010101010010",
						 "001010001001010101010000",
						 "001010001001010101001110",
						 "001010001001010101001100",
						 "001010001001010101001010",
						 "001010001001010101001000",
						 "001010001001010101000110",
						 "001010001001010101000100",
						 "001010001001010101000010",
						 "001010001001010101100000",
						 "001010001001010101011110",
						 "001010001001010101011100",
						 "001010001001010101011010",
						 "001010001001010101011000",
						 "001010001001010101010110",
						 "001010001001010101010100",
						 "001010001001010101010010",
						 "001010001001010101010000",
						 "001010001001010101001110",
						 "001010001001010101001100",
						 "001010001001010101001010",
						 "001010001001010101001000",
						 "001010001001010101000110",
						 "001010001001010101000100",
						 "001010001001010101000010",
						 "001010001001010101101111",
						 "001010001001010101101100",
						 "001010001001010101101001",
						 "001010001001010101100110",
						 "001010001001010101100011",
						 "001010001001010101100000",
						 "001010001001010101011101",
						 "001010001001010101011010",
						 "001010001001010101010111",
						 "001010001001010101010100",
						 "001010001001010101010001",
						 "001010001001010101001110",
						 "001010001001010101001011",
						 "001010001001010101001000",
						 "001010001001010101000101",
						 "001010001001010101000010",
						 "001010001001010101101111",
						 "001010001001010101101100",
						 "001010001001010101101001",
						 "001010001001010101100110",
						 "001010001001010101100011",
						 "001010001001010101100000",
						 "001010001001010101011101",
						 "001010001001010101011010",
						 "001010001001010101010111",
						 "001010001001010101010100",
						 "001010001001010101010001",
						 "001010001001010101001110",
						 "001010001001010101001011",
						 "001010001001010101001000",
						 "001010001001010101000101",
						 "001010001001010101000010",
						 "001010001001010101101111",
						 "001010001001010101101100",
						 "001010001001010101101001",
						 "001010001001010101100110",
						 "001010001001010101100011",
						 "001010001001010101100000",
						 "001010001001010101011101",
						 "001010001001010101011010",
						 "001010001001010101010111",
						 "001010001001010101010100",
						 "001010001001010101010001",
						 "001010001001010101001110",
						 "001010001001010101001011",
						 "001010001001010101001000",
						 "001010001001010101000101",
						 "001010001001010101000010",
						 "001010001001010101111110",
						 "001010001001010101111010",
						 "001010001001010101110110",
						 "001010001001010101110010",
						 "001010001001010101101110",
						 "001010001001010101101010",
						 "001010001001010101100110",
						 "001010001001010101100010",
						 "001010001001010101011110",
						 "001010001001010101011010",
						 "001010001001010101010110",
						 "001010001001010101010010",
						 "001010001001010101001110",
						 "001010001001010101001010",
						 "001010001001010101000110",
						 "001010001001010101000010",
						 "001010001001010101111110",
						 "001010001001010101111010",
						 "001010001001010101110110",
						 "001010001001010101110010",
						 "001010001001010101101110",
						 "001010001001010101101010",
						 "001010001001010101100110",
						 "001010001001010101100010",
						 "001010001001010101011110",
						 "001010001001010101011010",
						 "001010001001010101010110",
						 "001010001001010101010010",
						 "001010001001010101001110",
						 "001010001001010101001010",
						 "001010001001010101000110",
						 "001010001001010101000010",
						 "001010001001010101111110",
						 "001010001001010101111010",
						 "001010001001010101110110",
						 "001010001001010101110010",
						 "001010001001010101101110",
						 "001010001001010101101010",
						 "001010001001010101100110",
						 "001010001001010101100010",
						 "001010001001010101011110",
						 "001010001001010101011010",
						 "001010001001010101010110",
						 "001010001001010101010010",
						 "001010001001010101001110",
						 "001010001001010101001010",
						 "001010001001010101000110",
						 "001010001001010101000010",
						 "001010001001010110001101",
						 "001010001001010110001000",
						 "001010001001010110000011",
						 "001010001001010101111110",
						 "001010001001010101111001",
						 "001010001001010101110100",
						 "001010001001010101101111",
						 "001010001001010101101010",
						 "001010001001010101100101",
						 "001010001001010101100000",
						 "001010001001010101011011",
						 "001010001001010101010110",
						 "001010001001010101010001",
						 "001010001001010101001100",
						 "001010001001010101000111",
						 "001010001001010101000010",
						 "001010001001010110001101",
						 "001010001001010110001000",
						 "001010001001010110000011",
						 "001010001001010101111110",
						 "001010001001010101111001",
						 "001010001001010101110100",
						 "001010001001010101101111",
						 "001010001001010101101010",
						 "001010001001010101100101",
						 "001010001001010101100000",
						 "001010001001010101011011",
						 "001010001001010101010110",
						 "001010001001010101010001",
						 "001010001001010101001100",
						 "001010001001010101000111",
						 "001010001001010101000010",
						 "001010001001010110011100",
						 "001010001001010110010110",
						 "001010001001010110010000",
						 "001010001001010110001010",
						 "001010001001010110000100",
						 "001010001001010101111110",
						 "001010001001010101111000",
						 "001010001001010101110010",
						 "001010001001010101101100",
						 "001010001001010101100110",
						 "001010001001010101100000",
						 "001010001001010101011010",
						 "001010001001010101010100",
						 "001010001001010101001110",
						 "001010001001010101001000",
						 "001010001001010101000010",
						 "001010001001010110011100",
						 "001010001001010110010110",
						 "001010001001010110010000",
						 "001010001001010110001010",
						 "001010001001010110000100",
						 "001010001001010101111110",
						 "001010001001010101111000",
						 "001010001001010101110010",
						 "001010001001010101101100",
						 "001010001001010101100110",
						 "001010001001010101100000",
						 "001010001001010101011010",
						 "001010001001010101010100",
						 "001010001001010101001110",
						 "001010001001010101001000",
						 "001010001001010101000010",
						 "001010001001010110011100",
						 "001010001001010110010110",
						 "001010001001010110010000",
						 "001010001001010110001010",
						 "001010001001010110000100",
						 "001010001001010101111110",
						 "001010001001010101111000",
						 "001010001001010101110010",
						 "001010001001010101101100",
						 "001010001001010101100110",
						 "001010001001010101100000",
						 "001010001001010101011010",
						 "001010001001010101010100",
						 "001010001001010101001110",
						 "001010001001010101001000",
						 "001010001001010101000010",
						 "001010001001010110101011",
						 "001010001001010110100100",
						 "001010001001010110011101",
						 "001010001001010110010110",
						 "001010001001010110001111",
						 "001010001001010110001000",
						 "001010001001010110000001",
						 "001010001001010101111010",
						 "001010001001010101110011",
						 "001010001001010101101100",
						 "001010001001010101100101",
						 "001010001001010101011110",
						 "001010001001010101010111",
						 "001010001001010101010000",
						 "001010001001010101001001",
						 "001010001001010101000010",
						 "001010001001010110101011",
						 "001010001001010110100100",
						 "001010001001010110011101",
						 "001010001001010110010110",
						 "001010001001010110001111",
						 "001010001001010110001000",
						 "001010001001010110000001",
						 "001010001001010101111010",
						 "001010001001010101110011",
						 "001010001001010101101100",
						 "001010001001010101100101",
						 "001010001001010101011110",
						 "001010001001010101010111",
						 "001010001001010101010000",
						 "001010001001010101001001",
						 "001010001001010101000010",
						 "001010001001010110111010",
						 "001010001001010110110010",
						 "001010001001010110101010",
						 "001010001001010110100010",
						 "001010001001010110011010",
						 "001010001001010110010010",
						 "001010001001010110001010",
						 "001010001001010110000010",
						 "001010001001010101111010",
						 "001010001001010101110010",
						 "001010001001010101101010",
						 "001010001001010101100010",
						 "001010001001010101011010",
						 "001010001001010101010010",
						 "001010001001010101001010",
						 "001010001001010101000010",
						 "001010001001010110111010",
						 "001010001001010110110010",
						 "001010001001010110101010",
						 "001010001001010110100010",
						 "001010001001010110011010",
						 "001010001001010110010010",
						 "001010001001010110001010",
						 "001010001001010110000010",
						 "001010001001010101111010",
						 "001010001001010101110010",
						 "001010001001010101101010",
						 "001010001001010101100010",
						 "001010001001010101011010",
						 "001010001001010101010010",
						 "001010001001010101001010",
						 "001010001001010101000010",
						 "001010001001010110111010",
						 "001010001001010110110010",
						 "001010001001010110101010",
						 "001010001001010110100010",
						 "001010001001010110011010",
						 "001010001001010110010010",
						 "001010001001010110001010",
						 "001010001001010110000010",
						 "001010001001010101111010",
						 "001010001001010101110010",
						 "001010001001010101101010",
						 "001010001001010101100010",
						 "001010001001010101011010",
						 "001010001001010101010010",
						 "001010001001010101001010",
						 "001010001001010101000010",
						 "001010001001010111001001",
						 "001010001001010111000000",
						 "001010001001010110110111",
						 "001010001001010110101110",
						 "001010001001010110100101",
						 "001010001001010110011100",
						 "001010001001010110010011",
						 "001010001001010110001010",
						 "001010001001010110000001",
						 "001010001001010101111000",
						 "001010001001010101101111",
						 "001010001001010101100110",
						 "001010001001010101011101",
						 "001010001001010101010100",
						 "001010001001010101001011",
						 "001010001001010101000010",
						 "001010001001010111001001",
						 "001010001001010111000000",
						 "001010001001010110110111",
						 "001010001001010110101110",
						 "001010001001010110100101",
						 "001010001001010110011100",
						 "001010001001010110010011",
						 "001010001001010110001010",
						 "001010001001010110000001",
						 "001010001001010101111000",
						 "001010001001010101101111",
						 "001010001001010101100110",
						 "001010001001010101011101",
						 "001010001001010101010100",
						 "001010001001010101001011",
						 "001010001001010101000010",
						 "001010001001010111011000",
						 "001010001001010111001110",
						 "001010001001010111000100",
						 "001010001001010110111010",
						 "001010001001010110110000",
						 "001010001001010110100110",
						 "001010001001010110011100",
						 "001010001001010110010010",
						 "001010001001010110001000",
						 "001010001001010101111110",
						 "001010001001010101110100",
						 "001010001001010101101010",
						 "001010001001010101100000",
						 "001010001001010101010110",
						 "001010001001010101001100",
						 "001010001001010101000010",
						 "001010001001010111011000",
						 "001010001001010111001110",
						 "001010001001010111000100",
						 "001010001001010110111010",
						 "001010001001010110110000",
						 "001010001001010110100110",
						 "001010001001010110011100",
						 "001010001001010110010010",
						 "001010001001010110001000",
						 "001010001001010101111110",
						 "001010001001010101110100",
						 "001010001001010101101010",
						 "001010001001010101100000",
						 "001010001001010101010110",
						 "001010001001010101001100",
						 "001010001001010101000010",
						 "001010001001010111011000",
						 "001010001001010111001110",
						 "001010001001010111000100",
						 "001010001001010110111010",
						 "001010001001010110110000",
						 "001010001001010110100110",
						 "001010001001010110011100",
						 "001010001001010110010010",
						 "001010001001010110001000",
						 "001010001001010101111110",
						 "001010001001010101110100",
						 "001010001001010101101010",
						 "001010001001010101100000",
						 "001010001001010101010110",
						 "001010001001010101001100",
						 "001010001001010101000010",
						 "001010001001010111100111",
						 "001010001001010111011100",
						 "001010001001010111010001",
						 "001010001001010111000110",
						 "001010001001010110111011",
						 "001010001001010110110000",
						 "001010001001010110100101",
						 "001010001001010110011010",
						 "001010001001010110001111",
						 "001010001001010110000100",
						 "001010001001010101111001",
						 "001010001001010101101110",
						 "001010001001010101100011",
						 "001010001001010101011000",
						 "001010001001010101001101",
						 "001010001001010101000010",
						 "001010001001010111100111",
						 "001010001001010111011100",
						 "001010001001010111010001",
						 "001010001001010111000110",
						 "001010001001010110111011",
						 "001010001001010110110000",
						 "001010001001010110100101",
						 "001010001001010110011010",
						 "001010001001010110001111",
						 "001010001001010110000100",
						 "001010001001010101111001",
						 "001010001001010101101110",
						 "001010001001010101100011",
						 "001010001001010101011000",
						 "001010001001010101001101",
						 "001010001001010101000010",
						 "001010001001010111110110",
						 "001010001001010111101010",
						 "001010001001010111011110",
						 "001010001001010111010010",
						 "001010001001010111000110",
						 "001010001001010110111010",
						 "001010001001010110101110",
						 "001010001001010110100010",
						 "001010001001010110010110",
						 "001010001001010110001010",
						 "001010001001010101111110",
						 "001010001001010101110010",
						 "001010001001010101100110",
						 "001010001001010101011010",
						 "001010001001010101001110",
						 "001010001001010101000010",
						 "001010001001010111110110",
						 "001010001001010111101010",
						 "001010001001010111011110",
						 "001010001001010111010010",
						 "001010001001010111000110",
						 "001010001001010110111010",
						 "001010001001010110101110",
						 "001010001001010110100010",
						 "001010001001010110010110",
						 "001010001001010110001010",
						 "001010001001010101111110",
						 "001010001001010101110010",
						 "001010001001010101100110",
						 "001010001001010101011010",
						 "001010001001010101001110",
						 "001010001001010101000010",
						 "001010001001010111110110",
						 "001010001001010111101010",
						 "001010001001010111011110",
						 "001010001001010111010010",
						 "001010001001010111000110",
						 "001010001001010110111010",
						 "001010001001010110101110",
						 "001010001001010110100010",
						 "001010001001010110010110",
						 "001010001001010110001010",
						 "001010001001010101111110",
						 "001010001001010101110010",
						 "001010001001010101100110",
						 "001010001001010101011010",
						 "001010001001010101001110",
						 "001010001001010101000010",
						 "001010001001011000000101",
						 "001010001001010111111000",
						 "001010001001010111101011",
						 "001010001001010111011110",
						 "001010001001010111010001",
						 "001010001001010111000100",
						 "001010001001010110110111",
						 "001010001001010110101010",
						 "001010001001010110011101",
						 "001010001001010110010000",
						 "001010001001010110000011",
						 "001010001001010101110110",
						 "001010001001010101101001",
						 "001010001001010101011100",
						 "001010001001010101001111",
						 "001010001001010101000010",
						 "001010001001011000000101",
						 "001010001001010111111000",
						 "001010001001010111101011",
						 "001010001001010111011110",
						 "001010001001010111010001",
						 "001010001001010111000100",
						 "001010001001010110110111",
						 "001010001001010110101010",
						 "001010001001010110011101",
						 "001010001001010110010000",
						 "001010001001010110000011",
						 "001010001001010101110110",
						 "001010001001010101101001",
						 "001010001001010101011100",
						 "001010001001010101001111",
						 "001010001001010101000010",
						 "001010001001011000000101",
						 "001010001001010111111000",
						 "001010001001010111101011",
						 "001010001001010111011110",
						 "001010001001010111010001",
						 "001010001001010111000100",
						 "001010001001010110110111",
						 "001010001001010110101010",
						 "001010001001010110011101",
						 "001010001001010110010000",
						 "001010001001010110000011",
						 "001010001001010101110110",
						 "001010001001010101101001",
						 "001010001001010101011100",
						 "001010001001010101001111",
						 "001010001001010101000010",
						 "001010001001011000010100",
						 "001010001001011000000110",
						 "001010001001010111111000",
						 "001010001001010111101010",
						 "001010001001010111011100",
						 "001010001001010111001110",
						 "001010001001010111000000",
						 "001010001001010110110010",
						 "001010001001010110100100",
						 "001010001001010110010110",
						 "001010001001010110001000",
						 "001010001001010101111010",
						 "001010001001010101101100",
						 "001010001001010101011110",
						 "001010001001010101010000",
						 "001010001001010101000010",
						 "001010001001011000010100",
						 "001010001001011000000110",
						 "001010001001010111111000",
						 "001010001001010111101010",
						 "001010001001010111011100",
						 "001010001001010111001110",
						 "001010001001010111000000",
						 "001010001001010110110010",
						 "001010001001010110100100",
						 "001010001001010110010110",
						 "001010001001010110001000",
						 "001010001001010101111010",
						 "001010001001010101101100",
						 "001010001001010101011110",
						 "001010001001010101010000",
						 "001010001001010101000010",
						 "001010001001011000100011",
						 "001010001001011000010100",
						 "001010001001011000000101",
						 "001010001001010111110110",
						 "001010001001010111100111",
						 "001010001001010111011000",
						 "001010001001010111001001",
						 "001010001001010110111010",
						 "001010001001010110101011",
						 "001010001001010110011100",
						 "001010001001010110001101",
						 "001010001001010101111110",
						 "001010001001010101101111",
						 "001010001001010101100000",
						 "001010001001010101010001",
						 "001010001001010101000010",
						 "001010001001011000100011",
						 "001010001001011000010100",
						 "001010001001011000000101",
						 "001010001001010111110110",
						 "001010001001010111100111",
						 "001010001001010111011000",
						 "001010001001010111001001",
						 "001010001001010110111010",
						 "001010001001010110101011",
						 "001010001001010110011100",
						 "001010001001010110001101",
						 "001010001001010101111110",
						 "001010001001010101101111",
						 "001010001001010101100000",
						 "001010001001010101010001",
						 "001010001001010101000010",
						 "001010001001011000100011",
						 "001010001001011000010100",
						 "001010001001011000000101",
						 "001010001001010111110110",
						 "001010001001010111100111",
						 "001010001001010111011000",
						 "001010001001010111001001",
						 "001010001001010110111010",
						 "001010001001010110101011",
						 "001010001001010110011100",
						 "001010001001010110001101",
						 "001010001001010101111110",
						 "001010001001010101101111",
						 "001010001001010101100000",
						 "001010001001010101010001",
						 "001010001001010101000010",
						 "001010000110110101110100",
						 "001010000110110101100100",
						 "001010000110110101010100",
						 "001010000110110101000100",
						 "001010000110110100110100",
						 "001010000110110100100100",
						 "001010000110110100010100",
						 "001010000110110100000100",
						 "001010000110110011110100",
						 "001010000110110011100100",
						 "001010000110110011010100",
						 "001010000110110011000100",
						 "001010000110110010110100",
						 "001010000110110010100100",
						 "001010000110110010010100",
						 "001010000110110010000100",
						 "001010000110110101110100",
						 "001010000110110101100100",
						 "001010000110110101010100",
						 "001010000110110101000100",
						 "001010000110110100110100",
						 "001010000110110100100100",
						 "001010000110110100010100",
						 "001010000110110100000100",
						 "001010000110110011110100",
						 "001010000110110011100100",
						 "001010000110110011010100",
						 "001010000110110011000100",
						 "001010000110110010110100",
						 "001010000110110010100100",
						 "001010000110110010010100",
						 "001010000110110010000100",
						 "001010000110110110000011",
						 "001010000110110101110010",
						 "001010000110110101100001",
						 "001010000110110101010000",
						 "001010000110110100111111",
						 "001010000110110100101110",
						 "001010000110110100011101",
						 "001010000110110100001100",
						 "001010000110110011111011",
						 "001010000110110011101010",
						 "001010000110110011011001",
						 "001010000110110011001000",
						 "001010000110110010110111",
						 "001010000110110010100110",
						 "001010000110110010010101",
						 "001010000110110010000100",
						 "001010000110110110000011",
						 "001010000110110101110010",
						 "001010000110110101100001",
						 "001010000110110101010000",
						 "001010000110110100111111",
						 "001010000110110100101110",
						 "001010000110110100011101",
						 "001010000110110100001100",
						 "001010000110110011111011",
						 "001010000110110011101010",
						 "001010000110110011011001",
						 "001010000110110011001000",
						 "001010000110110010110111",
						 "001010000110110010100110",
						 "001010000110110010010101",
						 "001010000110110010000100",
						 "001010000110110110000011",
						 "001010000110110101110010",
						 "001010000110110101100001",
						 "001010000110110101010000",
						 "001010000110110100111111",
						 "001010000110110100101110",
						 "001010000110110100011101",
						 "001010000110110100001100",
						 "001010000110110011111011",
						 "001010000110110011101010",
						 "001010000110110011011001",
						 "001010000110110011001000",
						 "001010000110110010110111",
						 "001010000110110010100110",
						 "001010000110110010010101",
						 "001010000110110010000100",
						 "001010000110110110010010",
						 "001010000110110110000000",
						 "001010000110110101101110",
						 "001010000110110101011100",
						 "001010000110110101001010",
						 "001010000110110100111000",
						 "001010000110110100100110",
						 "001010000110110100010100",
						 "001010000110110100000010",
						 "001010000110110011110000",
						 "001010000110110011011110",
						 "001010000110110011001100",
						 "001010000110110010111010",
						 "001010000110110010101000",
						 "001010000110110010010110",
						 "001010000110110010000100",
						 "001010000110110110010010",
						 "001010000110110110000000",
						 "001010000110110101101110",
						 "001010000110110101011100",
						 "001010000110110101001010",
						 "001010000110110100111000",
						 "001010000110110100100110",
						 "001010000110110100010100",
						 "001010000110110100000010",
						 "001010000110110011110000",
						 "001010000110110011011110",
						 "001010000110110011001100",
						 "001010000110110010111010",
						 "001010000110110010101000",
						 "001010000110110010010110",
						 "001010000110110010000100",
						 "001010000110110110100001",
						 "001010000110110110001110",
						 "001010000110110101111011",
						 "001010000110110101101000",
						 "001010000110110101010101",
						 "001010000110110101000010",
						 "001010000110110100101111",
						 "001010000110110100011100",
						 "001010000110110100001001",
						 "001010000110110011110110",
						 "001010000110110011100011",
						 "001010000110110011010000",
						 "001010000110110010111101",
						 "001010000110110010101010",
						 "001010000110110010010111",
						 "001010000110110010000100",
						 "001010000110110110100001",
						 "001010000110110110001110",
						 "001010000110110101111011",
						 "001010000110110101101000",
						 "001010000110110101010101",
						 "001010000110110101000010",
						 "001010000110110100101111",
						 "001010000110110100011100",
						 "001010000110110100001001",
						 "001010000110110011110110",
						 "001010000110110011100011",
						 "001010000110110011010000",
						 "001010000110110010111101",
						 "001010000110110010101010",
						 "001010000110110010010111",
						 "001010000110110010000100",
						 "001010000110110110100001",
						 "001010000110110110001110",
						 "001010000110110101111011",
						 "001010000110110101101000",
						 "001010000110110101010101",
						 "001010000110110101000010",
						 "001010000110110100101111",
						 "001010000110110100011100",
						 "001010000110110100001001",
						 "001010000110110011110110",
						 "001010000110110011100011",
						 "001010000110110011010000",
						 "001010000110110010111101",
						 "001010000110110010101010",
						 "001010000110110010010111",
						 "001010000110110010000100",
						 "001010000110110110110000",
						 "001010000110110110011100",
						 "001010000110110110001000",
						 "001010000110110101110100",
						 "001010000110110101100000",
						 "001010000110110101001100",
						 "001010000110110100111000",
						 "001010000110110100100100",
						 "001010000110110100010000",
						 "001010000110110011111100",
						 "001010000110110011101000",
						 "001010000110110011010100",
						 "001010000110110011000000",
						 "001010000110110010101100",
						 "001010000110110010011000",
						 "001010000110110010000100",
						 "001010000110110110110000",
						 "001010000110110110011100",
						 "001010000110110110001000",
						 "001010000110110101110100",
						 "001010000110110101100000",
						 "001010000110110101001100",
						 "001010000110110100111000",
						 "001010000110110100100100",
						 "001010000110110100010000",
						 "001010000110110011111100",
						 "001010000110110011101000",
						 "001010000110110011010100",
						 "001010000110110011000000",
						 "001010000110110010101100",
						 "001010000110110010011000",
						 "001010000110110010000100",
						 "001010000110110110111111",
						 "001010000110110110101010",
						 "001010000110110110010101",
						 "001010000110110110000000",
						 "001010000110110101101011",
						 "001010000110110101010110",
						 "001010000110110101000001",
						 "001010000110110100101100",
						 "001010000110110100010111",
						 "001010000110110100000010",
						 "001010000110110011101101",
						 "001010000110110011011000",
						 "001010000110110011000011",
						 "001010000110110010101110",
						 "001010000110110010011001",
						 "001010000110110010000100",
						 "001010000110110110111111",
						 "001010000110110110101010",
						 "001010000110110110010101",
						 "001010000110110110000000",
						 "001010000110110101101011",
						 "001010000110110101010110",
						 "001010000110110101000001",
						 "001010000110110100101100",
						 "001010000110110100010111",
						 "001010000110110100000010",
						 "001010000110110011101101",
						 "001010000110110011011000",
						 "001010000110110011000011",
						 "001010000110110010101110",
						 "001010000110110010011001",
						 "001010000110110010000100",
						 "001010000110110110111111",
						 "001010000110110110101010",
						 "001010000110110110010101",
						 "001010000110110110000000",
						 "001010000110110101101011",
						 "001010000110110101010110",
						 "001010000110110101000001",
						 "001010000110110100101100",
						 "001010000110110100010111",
						 "001010000110110100000010",
						 "001010000110110011101101",
						 "001010000110110011011000",
						 "001010000110110011000011",
						 "001010000110110010101110",
						 "001010000110110010011001",
						 "001010000110110010000100",
						 "001010000110110111001110",
						 "001010000110110110111000",
						 "001010000110110110100010",
						 "001010000110110110001100",
						 "001010000110110101110110",
						 "001010000110110101100000",
						 "001010000110110101001010",
						 "001010000110110100110100",
						 "001010000110110100011110",
						 "001010000110110100001000",
						 "001010000110110011110010",
						 "001010000110110011011100",
						 "001010000110110011000110",
						 "001010000110110010110000",
						 "001010000110110010011010",
						 "001010000110110010000100",
						 "001010000110110111001110",
						 "001010000110110110111000",
						 "001010000110110110100010",
						 "001010000110110110001100",
						 "001010000110110101110110",
						 "001010000110110101100000",
						 "001010000110110101001010",
						 "001010000110110100110100",
						 "001010000110110100011110",
						 "001010000110110100001000",
						 "001010000110110011110010",
						 "001010000110110011011100",
						 "001010000110110011000110",
						 "001010000110110010110000",
						 "001010000110110010011010",
						 "001010000110110010000100",
						 "001010000110110111001110",
						 "001010000110110110111000",
						 "001010000110110110100010",
						 "001010000110110110001100",
						 "001010000110110101110110",
						 "001010000110110101100000",
						 "001010000110110101001010",
						 "001010000110110100110100",
						 "001010000110110100011110",
						 "001010000110110100001000",
						 "001010000110110011110010",
						 "001010000110110011011100",
						 "001010000110110011000110",
						 "001010000110110010110000",
						 "001010000110110010011010",
						 "001010000110110010000100",
						 "001010000110110111011101",
						 "001010000110110111000110",
						 "001010000110110110101111",
						 "001010000110110110011000",
						 "001010000110110110000001",
						 "001010000110110101101010",
						 "001010000110110101010011",
						 "001010000110110100111100",
						 "001010000110110100100101",
						 "001010000110110100001110",
						 "001010000110110011110111",
						 "001010000110110011100000",
						 "001010000110110011001001",
						 "001010000110110010110010",
						 "001010000110110010011011",
						 "001010000110110010000100",
						 "001010000110110111011101",
						 "001010000110110111000110",
						 "001010000110110110101111",
						 "001010000110110110011000",
						 "001010000110110110000001",
						 "001010000110110101101010",
						 "001010000110110101010011",
						 "001010000110110100111100",
						 "001010000110110100100101",
						 "001010000110110100001110",
						 "001010000110110011110111",
						 "001010000110110011100000",
						 "001010000110110011001001",
						 "001010000110110010110010",
						 "001010000110110010011011",
						 "001010000110110010000100",
						 "001010000110110111101100",
						 "001010000110110111010100",
						 "001010000110110110111100",
						 "001010000110110110100100",
						 "001010000110110110001100",
						 "001010000110110101110100",
						 "001010000110110101011100",
						 "001010000110110101000100",
						 "001010000110110100101100",
						 "001010000110110100010100",
						 "001010000110110011111100",
						 "001010000110110011100100",
						 "001010000110110011001100",
						 "001010000110110010110100",
						 "001010000110110010011100",
						 "001010000110110010000100",
						 "001010000110110111101100",
						 "001010000110110111010100",
						 "001010000110110110111100",
						 "001010000110110110100100",
						 "001010000110110110001100",
						 "001010000110110101110100",
						 "001010000110110101011100",
						 "001010000110110101000100",
						 "001010000110110100101100",
						 "001010000110110100010100",
						 "001010000110110011111100",
						 "001010000110110011100100",
						 "001010000110110011001100",
						 "001010000110110010110100",
						 "001010000110110010011100",
						 "001010000110110010000100",
						 "001010000110110111101100",
						 "001010000110110111010100",
						 "001010000110110110111100",
						 "001010000110110110100100",
						 "001010000110110110001100",
						 "001010000110110101110100",
						 "001010000110110101011100",
						 "001010000110110101000100",
						 "001010000110110100101100",
						 "001010000110110100010100",
						 "001010000110110011111100",
						 "001010000110110011100100",
						 "001010000110110011001100",
						 "001010000110110010110100",
						 "001010000110110010011100",
						 "001010000110110010000100",
						 "001010000110110111111011",
						 "001010000110110111100010",
						 "001010000110110111001001",
						 "001010000110110110110000",
						 "001010000110110110010111",
						 "001010000110110101111110",
						 "001010000110110101100101",
						 "001010000110110101001100",
						 "001010000110110100110011",
						 "001010000110110100011010",
						 "001010000110110100000001",
						 "001010000110110011101000",
						 "001010000110110011001111",
						 "001010000110110010110110",
						 "001010000110110010011101",
						 "001010000110110010000100",
						 "001010000110110111111011",
						 "001010000110110111100010",
						 "001010000110110111001001",
						 "001010000110110110110000",
						 "001010000110110110010111",
						 "001010000110110101111110",
						 "001010000110110101100101",
						 "001010000110110101001100",
						 "001010000110110100110011",
						 "001010000110110100011010",
						 "001010000110110100000001",
						 "001010000110110011101000",
						 "001010000110110011001111",
						 "001010000110110010110110",
						 "001010000110110010011101",
						 "001010000110110010000100",
						 "001010000110111000001010",
						 "001010000110110111110000",
						 "001010000110110111010110",
						 "001010000110110110111100",
						 "001010000110110110100010",
						 "001010000110110110001000",
						 "001010000110110101101110",
						 "001010000110110101010100",
						 "001010000110110100111010",
						 "001010000110110100100000",
						 "001010000110110100000110",
						 "001010000110110011101100",
						 "001010000110110011010010",
						 "001010000110110010111000",
						 "001010000110110010011110",
						 "001010000110110010000100",
						 "001010000110111000001010",
						 "001010000110110111110000",
						 "001010000110110111010110",
						 "001010000110110110111100",
						 "001010000110110110100010",
						 "001010000110110110001000",
						 "001010000110110101101110",
						 "001010000110110101010100",
						 "001010000110110100111010",
						 "001010000110110100100000",
						 "001010000110110100000110",
						 "001010000110110011101100",
						 "001010000110110011010010",
						 "001010000110110010111000",
						 "001010000110110010011110",
						 "001010000110110010000100",
						 "001010000110111000001010",
						 "001010000110110111110000",
						 "001010000110110111010110",
						 "001010000110110110111100",
						 "001010000110110110100010",
						 "001010000110110110001000",
						 "001010000110110101101110",
						 "001010000110110101010100",
						 "001010000110110100111010",
						 "001010000110110100100000",
						 "001010000110110100000110",
						 "001010000110110011101100",
						 "001010000110110011010010",
						 "001010000110110010111000",
						 "001010000110110010011110",
						 "001010000110110010000100",
						 "001010000110111000011001",
						 "001010000110110111111110",
						 "001010000110110111100011",
						 "001010000110110111001000",
						 "001010000110110110101101",
						 "001010000110110110010010",
						 "001010000110110101110111",
						 "001010000110110101011100",
						 "001010000110110101000001",
						 "001010000110110100100110",
						 "001010000110110100001011",
						 "001010000110110011110000",
						 "001010000110110011010101",
						 "001010000110110010111010",
						 "001010000110110010011111",
						 "001010000110110010000100",
						 "001010000110111000011001",
						 "001010000110110111111110",
						 "001010000110110111100011",
						 "001010000110110111001000",
						 "001010000110110110101101",
						 "001010000110110110010010",
						 "001010000110110101110111",
						 "001010000110110101011100",
						 "001010000110110101000001",
						 "001010000110110100100110",
						 "001010000110110100001011",
						 "001010000110110011110000",
						 "001010000110110011010101",
						 "001010000110110010111010",
						 "001010000110110010011111",
						 "001010000110110010000100",
						 "001010000100010101101010",
						 "001010000100010101001110",
						 "001010000100010100110010",
						 "001010000100010100010110",
						 "001010000100010011111010",
						 "001010000100010011011110",
						 "001010000100010011000010",
						 "001010000100010010100110",
						 "001010000100010010001010",
						 "001010000100010001101110",
						 "001010000100010001010010",
						 "001010000100010000110110",
						 "001010000100010000011010",
						 "001010000100001111111110",
						 "001010000100001111100010",
						 "001010000100001111000110",
						 "001010000100010101101010",
						 "001010000100010101001110",
						 "001010000100010100110010",
						 "001010000100010100010110",
						 "001010000100010011111010",
						 "001010000100010011011110",
						 "001010000100010011000010",
						 "001010000100010010100110",
						 "001010000100010010001010",
						 "001010000100010001101110",
						 "001010000100010001010010",
						 "001010000100010000110110",
						 "001010000100010000011010",
						 "001010000100001111111110",
						 "001010000100001111100010",
						 "001010000100001111000110",
						 "001010000100010101101010",
						 "001010000100010101001110",
						 "001010000100010100110010",
						 "001010000100010100010110",
						 "001010000100010011111010",
						 "001010000100010011011110",
						 "001010000100010011000010",
						 "001010000100010010100110",
						 "001010000100010010001010",
						 "001010000100010001101110",
						 "001010000100010001010010",
						 "001010000100010000110110",
						 "001010000100010000011010",
						 "001010000100001111111110",
						 "001010000100001111100010",
						 "001010000100001111000110",
						 "001010000100010101111001",
						 "001010000100010101011100",
						 "001010000100010100111111",
						 "001010000100010100100010",
						 "001010000100010100000101",
						 "001010000100010011101000",
						 "001010000100010011001011",
						 "001010000100010010101110",
						 "001010000100010010010001",
						 "001010000100010001110100",
						 "001010000100010001010111",
						 "001010000100010000111010",
						 "001010000100010000011101",
						 "001010000100010000000000",
						 "001010000100001111100011",
						 "001010000100001111000110",
						 "001010000100010101111001",
						 "001010000100010101011100",
						 "001010000100010100111111",
						 "001010000100010100100010",
						 "001010000100010100000101",
						 "001010000100010011101000",
						 "001010000100010011001011",
						 "001010000100010010101110",
						 "001010000100010010010001",
						 "001010000100010001110100",
						 "001010000100010001010111",
						 "001010000100010000111010",
						 "001010000100010000011101",
						 "001010000100010000000000",
						 "001010000100001111100011",
						 "001010000100001111000110",
						 "001010000100010101111001",
						 "001010000100010101011100",
						 "001010000100010100111111",
						 "001010000100010100100010",
						 "001010000100010100000101",
						 "001010000100010011101000",
						 "001010000100010011001011",
						 "001010000100010010101110",
						 "001010000100010010010001",
						 "001010000100010001110100",
						 "001010000100010001010111",
						 "001010000100010000111010",
						 "001010000100010000011101",
						 "001010000100010000000000",
						 "001010000100001111100011",
						 "001010000100001111000110",
						 "001010000100010110001000",
						 "001010000100010101101010",
						 "001010000100010101001100",
						 "001010000100010100101110",
						 "001010000100010100010000",
						 "001010000100010011110010",
						 "001010000100010011010100",
						 "001010000100010010110110",
						 "001010000100010010011000",
						 "001010000100010001111010",
						 "001010000100010001011100",
						 "001010000100010000111110",
						 "001010000100010000100000",
						 "001010000100010000000010",
						 "001010000100001111100100",
						 "001010000100001111000110",
						 "001010000100010110001000",
						 "001010000100010101101010",
						 "001010000100010101001100",
						 "001010000100010100101110",
						 "001010000100010100010000",
						 "001010000100010011110010",
						 "001010000100010011010100",
						 "001010000100010010110110",
						 "001010000100010010011000",
						 "001010000100010001111010",
						 "001010000100010001011100",
						 "001010000100010000111110",
						 "001010000100010000100000",
						 "001010000100010000000010",
						 "001010000100001111100100",
						 "001010000100001111000110",
						 "001010000100010110010111",
						 "001010000100010101111000",
						 "001010000100010101011001",
						 "001010000100010100111010",
						 "001010000100010100011011",
						 "001010000100010011111100",
						 "001010000100010011011101",
						 "001010000100010010111110",
						 "001010000100010010011111",
						 "001010000100010010000000",
						 "001010000100010001100001",
						 "001010000100010001000010",
						 "001010000100010000100011",
						 "001010000100010000000100",
						 "001010000100001111100101",
						 "001010000100001111000110",
						 "001010000100010110010111",
						 "001010000100010101111000",
						 "001010000100010101011001",
						 "001010000100010100111010",
						 "001010000100010100011011",
						 "001010000100010011111100",
						 "001010000100010011011101",
						 "001010000100010010111110",
						 "001010000100010010011111",
						 "001010000100010010000000",
						 "001010000100010001100001",
						 "001010000100010001000010",
						 "001010000100010000100011",
						 "001010000100010000000100",
						 "001010000100001111100101",
						 "001010000100001111000110",
						 "001010000100010110010111",
						 "001010000100010101111000",
						 "001010000100010101011001",
						 "001010000100010100111010",
						 "001010000100010100011011",
						 "001010000100010011111100",
						 "001010000100010011011101",
						 "001010000100010010111110",
						 "001010000100010010011111",
						 "001010000100010010000000",
						 "001010000100010001100001",
						 "001010000100010001000010",
						 "001010000100010000100011",
						 "001010000100010000000100",
						 "001010000100001111100101",
						 "001010000100001111000110",
						 "001010000100010110100110",
						 "001010000100010110000110",
						 "001010000100010101100110",
						 "001010000100010101000110",
						 "001010000100010100100110",
						 "001010000100010100000110",
						 "001010000100010011100110",
						 "001010000100010011000110",
						 "001010000100010010100110",
						 "001010000100010010000110",
						 "001010000100010001100110",
						 "001010000100010001000110",
						 "001010000100010000100110",
						 "001010000100010000000110",
						 "001010000100001111100110",
						 "001010000100001111000110",
						 "001010000100010110100110",
						 "001010000100010110000110",
						 "001010000100010101100110",
						 "001010000100010101000110",
						 "001010000100010100100110",
						 "001010000100010100000110",
						 "001010000100010011100110",
						 "001010000100010011000110",
						 "001010000100010010100110",
						 "001010000100010010000110",
						 "001010000100010001100110",
						 "001010000100010001000110",
						 "001010000100010000100110",
						 "001010000100010000000110",
						 "001010000100001111100110",
						 "001010000100001111000110",
						 "001010000100010110110101",
						 "001010000100010110010100",
						 "001010000100010101110011",
						 "001010000100010101010010",
						 "001010000100010100110001",
						 "001010000100010100010000",
						 "001010000100010011101111",
						 "001010000100010011001110",
						 "001010000100010010101101",
						 "001010000100010010001100",
						 "001010000100010001101011",
						 "001010000100010001001010",
						 "001010000100010000101001",
						 "001010000100010000001000",
						 "001010000100001111100111",
						 "001010000100001111000110",
						 "001010000100010110110101",
						 "001010000100010110010100",
						 "001010000100010101110011",
						 "001010000100010101010010",
						 "001010000100010100110001",
						 "001010000100010100010000",
						 "001010000100010011101111",
						 "001010000100010011001110",
						 "001010000100010010101101",
						 "001010000100010010001100",
						 "001010000100010001101011",
						 "001010000100010001001010",
						 "001010000100010000101001",
						 "001010000100010000001000",
						 "001010000100001111100111",
						 "001010000100001111000110",
						 "001010000100010110110101",
						 "001010000100010110010100",
						 "001010000100010101110011",
						 "001010000100010101010010",
						 "001010000100010100110001",
						 "001010000100010100010000",
						 "001010000100010011101111",
						 "001010000100010011001110",
						 "001010000100010010101101",
						 "001010000100010010001100",
						 "001010000100010001101011",
						 "001010000100010001001010",
						 "001010000100010000101001",
						 "001010000100010000001000",
						 "001010000100001111100111",
						 "001010000100001111000110",
						 "001010000100010111000100",
						 "001010000100010110100010",
						 "001010000100010110000000",
						 "001010000100010101011110",
						 "001010000100010100111100",
						 "001010000100010100011010",
						 "001010000100010011111000",
						 "001010000100010011010110",
						 "001010000100010010110100",
						 "001010000100010010010010",
						 "001010000100010001110000",
						 "001010000100010001001110",
						 "001010000100010000101100",
						 "001010000100010000001010",
						 "001010000100001111101000",
						 "001010000100001111000110",
						 "001010000100010111000100",
						 "001010000100010110100010",
						 "001010000100010110000000",
						 "001010000100010101011110",
						 "001010000100010100111100",
						 "001010000100010100011010",
						 "001010000100010011111000",
						 "001010000100010011010110",
						 "001010000100010010110100",
						 "001010000100010010010010",
						 "001010000100010001110000",
						 "001010000100010001001110",
						 "001010000100010000101100",
						 "001010000100010000001010",
						 "001010000100001111101000",
						 "001010000100001111000110",
						 "001010000100010111010011",
						 "001010000100010110110000",
						 "001010000100010110001101",
						 "001010000100010101101010",
						 "001010000100010101000111",
						 "001010000100010100100100",
						 "001010000100010100000001",
						 "001010000100010011011110",
						 "001010000100010010111011",
						 "001010000100010010011000",
						 "001010000100010001110101",
						 "001010000100010001010010",
						 "001010000100010000101111",
						 "001010000100010000001100",
						 "001010000100001111101001",
						 "001010000100001111000110",
						 "001010000100010111010011",
						 "001010000100010110110000",
						 "001010000100010110001101",
						 "001010000100010101101010",
						 "001010000100010101000111",
						 "001010000100010100100100",
						 "001010000100010100000001",
						 "001010000100010011011110",
						 "001010000100010010111011",
						 "001010000100010010011000",
						 "001010000100010001110101",
						 "001010000100010001010010",
						 "001010000100010000101111",
						 "001010000100010000001100",
						 "001010000100001111101001",
						 "001010000100001111000110",
						 "001010000100010111010011",
						 "001010000100010110110000",
						 "001010000100010110001101",
						 "001010000100010101101010",
						 "001010000100010101000111",
						 "001010000100010100100100",
						 "001010000100010100000001",
						 "001010000100010011011110",
						 "001010000100010010111011",
						 "001010000100010010011000",
						 "001010000100010001110101",
						 "001010000100010001010010",
						 "001010000100010000101111",
						 "001010000100010000001100",
						 "001010000100001111101001",
						 "001010000100001111000110",
						 "001010000001110100100100",
						 "001010000001110100000000",
						 "001010000001110011011100",
						 "001010000001110010111000",
						 "001010000001110010010100",
						 "001010000001110001110000",
						 "001010000001110001001100",
						 "001010000001110000101000",
						 "001010000001110000000100",
						 "001010000001101111100000",
						 "001010000001101110111100",
						 "001010000001101110011000",
						 "001010000001101101110100",
						 "001010000001101101010000",
						 "001010000001101100101100",
						 "001010000001101100001000",
						 "001010000001110100100100",
						 "001010000001110100000000",
						 "001010000001110011011100",
						 "001010000001110010111000",
						 "001010000001110010010100",
						 "001010000001110001110000",
						 "001010000001110001001100",
						 "001010000001110000101000",
						 "001010000001110000000100",
						 "001010000001101111100000",
						 "001010000001101110111100",
						 "001010000001101110011000",
						 "001010000001101101110100",
						 "001010000001101101010000",
						 "001010000001101100101100",
						 "001010000001101100001000",
						 "001010000001110100100100",
						 "001010000001110100000000",
						 "001010000001110011011100",
						 "001010000001110010111000",
						 "001010000001110010010100",
						 "001010000001110001110000",
						 "001010000001110001001100",
						 "001010000001110000101000",
						 "001010000001110000000100",
						 "001010000001101111100000",
						 "001010000001101110111100",
						 "001010000001101110011000",
						 "001010000001101101110100",
						 "001010000001101101010000",
						 "001010000001101100101100",
						 "001010000001101100001000",
						 "001010000001110100110011",
						 "001010000001110100001110",
						 "001010000001110011101001",
						 "001010000001110011000100",
						 "001010000001110010011111",
						 "001010000001110001111010",
						 "001010000001110001010101",
						 "001010000001110000110000",
						 "001010000001110000001011",
						 "001010000001101111100110",
						 "001010000001101111000001",
						 "001010000001101110011100",
						 "001010000001101101110111",
						 "001010000001101101010010",
						 "001010000001101100101101",
						 "001010000001101100001000",
						 "001010000001110100110011",
						 "001010000001110100001110",
						 "001010000001110011101001",
						 "001010000001110011000100",
						 "001010000001110010011111",
						 "001010000001110001111010",
						 "001010000001110001010101",
						 "001010000001110000110000",
						 "001010000001110000001011",
						 "001010000001101111100110",
						 "001010000001101111000001",
						 "001010000001101110011100",
						 "001010000001101101110111",
						 "001010000001101101010010",
						 "001010000001101100101101",
						 "001010000001101100001000",
						 "001010000001110101000010",
						 "001010000001110100011100",
						 "001010000001110011110110",
						 "001010000001110011010000",
						 "001010000001110010101010",
						 "001010000001110010000100",
						 "001010000001110001011110",
						 "001010000001110000111000",
						 "001010000001110000010010",
						 "001010000001101111101100",
						 "001010000001101111000110",
						 "001010000001101110100000",
						 "001010000001101101111010",
						 "001010000001101101010100",
						 "001010000001101100101110",
						 "001010000001101100001000",
						 "001010000001110101000010",
						 "001010000001110100011100",
						 "001010000001110011110110",
						 "001010000001110011010000",
						 "001010000001110010101010",
						 "001010000001110010000100",
						 "001010000001110001011110",
						 "001010000001110000111000",
						 "001010000001110000010010",
						 "001010000001101111101100",
						 "001010000001101111000110",
						 "001010000001101110100000",
						 "001010000001101101111010",
						 "001010000001101101010100",
						 "001010000001101100101110",
						 "001010000001101100001000",
						 "001010000001110101000010",
						 "001010000001110100011100",
						 "001010000001110011110110",
						 "001010000001110011010000",
						 "001010000001110010101010",
						 "001010000001110010000100",
						 "001010000001110001011110",
						 "001010000001110000111000",
						 "001010000001110000010010",
						 "001010000001101111101100",
						 "001010000001101111000110",
						 "001010000001101110100000",
						 "001010000001101101111010",
						 "001010000001101101010100",
						 "001010000001101100101110",
						 "001010000001101100001000",
						 "001010000001110101010001",
						 "001010000001110100101010",
						 "001010000001110100000011",
						 "001010000001110011011100",
						 "001010000001110010110101",
						 "001010000001110010001110",
						 "001010000001110001100111",
						 "001010000001110001000000",
						 "001010000001110000011001",
						 "001010000001101111110010",
						 "001010000001101111001011",
						 "001010000001101110100100",
						 "001010000001101101111101",
						 "001010000001101101010110",
						 "001010000001101100101111",
						 "001010000001101100001000",
						 "001010000001110101010001",
						 "001010000001110100101010",
						 "001010000001110100000011",
						 "001010000001110011011100",
						 "001010000001110010110101",
						 "001010000001110010001110",
						 "001010000001110001100111",
						 "001010000001110001000000",
						 "001010000001110000011001",
						 "001010000001101111110010",
						 "001010000001101111001011",
						 "001010000001101110100100",
						 "001010000001101101111101",
						 "001010000001101101010110",
						 "001010000001101100101111",
						 "001010000001101100001000",
						 "001010000001110101100000",
						 "001010000001110100111000",
						 "001010000001110100010000",
						 "001010000001110011101000",
						 "001010000001110011000000",
						 "001010000001110010011000",
						 "001010000001110001110000",
						 "001010000001110001001000",
						 "001010000001110000100000",
						 "001010000001101111111000",
						 "001010000001101111010000",
						 "001010000001101110101000",
						 "001010000001101110000000",
						 "001010000001101101011000",
						 "001010000001101100110000",
						 "001010000001101100001000",
						 "001010000001110101100000",
						 "001010000001110100111000",
						 "001010000001110100010000",
						 "001010000001110011101000",
						 "001010000001110011000000",
						 "001010000001110010011000",
						 "001010000001110001110000",
						 "001010000001110001001000",
						 "001010000001110000100000",
						 "001010000001101111111000",
						 "001010000001101111010000",
						 "001010000001101110101000",
						 "001010000001101110000000",
						 "001010000001101101011000",
						 "001010000001101100110000",
						 "001010000001101100001000",
						 "001010000001110101100000",
						 "001010000001110100111000",
						 "001010000001110100010000",
						 "001010000001110011101000",
						 "001010000001110011000000",
						 "001010000001110010011000",
						 "001010000001110001110000",
						 "001010000001110001001000",
						 "001010000001110000100000",
						 "001010000001101111111000",
						 "001010000001101111010000",
						 "001010000001101110101000",
						 "001010000001101110000000",
						 "001010000001101101011000",
						 "001010000001101100110000",
						 "001010000001101100001000",
						 "001010000001110101101111",
						 "001010000001110101000110",
						 "001010000001110100011101",
						 "001010000001110011110100",
						 "001010000001110011001011",
						 "001010000001110010100010",
						 "001010000001110001111001",
						 "001010000001110001010000",
						 "001010000001110000100111",
						 "001010000001101111111110",
						 "001010000001101111010101",
						 "001010000001101110101100",
						 "001010000001101110000011",
						 "001010000001101101011010",
						 "001010000001101100110001",
						 "001010000001101100001000",
						 "001010000001110101101111",
						 "001010000001110101000110",
						 "001010000001110100011101",
						 "001010000001110011110100",
						 "001010000001110011001011",
						 "001010000001110010100010",
						 "001010000001110001111001",
						 "001010000001110001010000",
						 "001010000001110000100111",
						 "001010000001101111111110",
						 "001010000001101111010101",
						 "001010000001101110101100",
						 "001010000001101110000011",
						 "001010000001101101011010",
						 "001010000001101100110001",
						 "001010000001101100001000",
						 "001010000001110101101111",
						 "001010000001110101000110",
						 "001010000001110100011101",
						 "001010000001110011110100",
						 "001010000001110011001011",
						 "001010000001110010100010",
						 "001010000001110001111001",
						 "001010000001110001010000",
						 "001010000001110000100111",
						 "001010000001101111111110",
						 "001010000001101111010101",
						 "001010000001101110101100",
						 "001010000001101110000011",
						 "001010000001101101011010",
						 "001010000001101100110001",
						 "001010000001101100001000",
						 "001010000001110101111110",
						 "001010000001110101010100",
						 "001010000001110100101010",
						 "001010000001110100000000",
						 "001010000001110011010110",
						 "001010000001110010101100",
						 "001010000001110010000010",
						 "001010000001110001011000",
						 "001010000001110000101110",
						 "001010000001110000000100",
						 "001010000001101111011010",
						 "001010000001101110110000",
						 "001010000001101110000110",
						 "001010000001101101011100",
						 "001010000001101100110010",
						 "001010000001101100001000",
						 "001001111111010011000000",
						 "001001111111010010010110",
						 "001001111111010001101100",
						 "001001111111010001000010",
						 "001001111111010000011000",
						 "001001111111001111101110",
						 "001001111111001111000100",
						 "001001111111001110011010",
						 "001001111111001101110000",
						 "001001111111001101000110",
						 "001001111111001100011100",
						 "001001111111001011110010",
						 "001001111111001011001000",
						 "001001111111001010011110",
						 "001001111111001001110100",
						 "001001111111001001001010",
						 "001001111111010011001111",
						 "001001111111010010100100",
						 "001001111111010001111001",
						 "001001111111010001001110",
						 "001001111111010000100011",
						 "001001111111001111111000",
						 "001001111111001111001101",
						 "001001111111001110100010",
						 "001001111111001101110111",
						 "001001111111001101001100",
						 "001001111111001100100001",
						 "001001111111001011110110",
						 "001001111111001011001011",
						 "001001111111001010100000",
						 "001001111111001001110101",
						 "001001111111001001001010",
						 "001001111111010011001111",
						 "001001111111010010100100",
						 "001001111111010001111001",
						 "001001111111010001001110",
						 "001001111111010000100011",
						 "001001111111001111111000",
						 "001001111111001111001101",
						 "001001111111001110100010",
						 "001001111111001101110111",
						 "001001111111001101001100",
						 "001001111111001100100001",
						 "001001111111001011110110",
						 "001001111111001011001011",
						 "001001111111001010100000",
						 "001001111111001001110101",
						 "001001111111001001001010",
						 "001001111111010011001111",
						 "001001111111010010100100",
						 "001001111111010001111001",
						 "001001111111010001001110",
						 "001001111111010000100011",
						 "001001111111001111111000",
						 "001001111111001111001101",
						 "001001111111001110100010",
						 "001001111111001101110111",
						 "001001111111001101001100",
						 "001001111111001100100001",
						 "001001111111001011110110",
						 "001001111111001011001011",
						 "001001111111001010100000",
						 "001001111111001001110101",
						 "001001111111001001001010",
						 "001001111111010011011110",
						 "001001111111010010110010",
						 "001001111111010010000110",
						 "001001111111010001011010",
						 "001001111111010000101110",
						 "001001111111010000000010",
						 "001001111111001111010110",
						 "001001111111001110101010",
						 "001001111111001101111110",
						 "001001111111001101010010",
						 "001001111111001100100110",
						 "001001111111001011111010",
						 "001001111111001011001110",
						 "001001111111001010100010",
						 "001001111111001001110110",
						 "001001111111001001001010",
						 "001001111111010011011110",
						 "001001111111010010110010",
						 "001001111111010010000110",
						 "001001111111010001011010",
						 "001001111111010000101110",
						 "001001111111010000000010",
						 "001001111111001111010110",
						 "001001111111001110101010",
						 "001001111111001101111110",
						 "001001111111001101010010",
						 "001001111111001100100110",
						 "001001111111001011111010",
						 "001001111111001011001110",
						 "001001111111001010100010",
						 "001001111111001001110110",
						 "001001111111001001001010",
						 "001001111111010011101101",
						 "001001111111010011000000",
						 "001001111111010010010011",
						 "001001111111010001100110",
						 "001001111111010000111001",
						 "001001111111010000001100",
						 "001001111111001111011111",
						 "001001111111001110110010",
						 "001001111111001110000101",
						 "001001111111001101011000",
						 "001001111111001100101011",
						 "001001111111001011111110",
						 "001001111111001011010001",
						 "001001111111001010100100",
						 "001001111111001001110111",
						 "001001111111001001001010",
						 "001001111111010011101101",
						 "001001111111010011000000",
						 "001001111111010010010011",
						 "001001111111010001100110",
						 "001001111111010000111001",
						 "001001111111010000001100",
						 "001001111111001111011111",
						 "001001111111001110110010",
						 "001001111111001110000101",
						 "001001111111001101011000",
						 "001001111111001100101011",
						 "001001111111001011111110",
						 "001001111111001011010001",
						 "001001111111001010100100",
						 "001001111111001001110111",
						 "001001111111001001001010",
						 "001001111111010011101101",
						 "001001111111010011000000",
						 "001001111111010010010011",
						 "001001111111010001100110",
						 "001001111111010000111001",
						 "001001111111010000001100",
						 "001001111111001111011111",
						 "001001111111001110110010",
						 "001001111111001110000101",
						 "001001111111001101011000",
						 "001001111111001100101011",
						 "001001111111001011111110",
						 "001001111111001011010001",
						 "001001111111001010100100",
						 "001001111111001001110111",
						 "001001111111001001001010",
						 "001001111111010011111100",
						 "001001111111010011001110",
						 "001001111111010010100000",
						 "001001111111010001110010",
						 "001001111111010001000100",
						 "001001111111010000010110",
						 "001001111111001111101000",
						 "001001111111001110111010",
						 "001001111111001110001100",
						 "001001111111001101011110",
						 "001001111111001100110000",
						 "001001111111001100000010",
						 "001001111111001011010100",
						 "001001111111001010100110",
						 "001001111111001001111000",
						 "001001111111001001001010",
						 "001001111111010011111100",
						 "001001111111010011001110",
						 "001001111111010010100000",
						 "001001111111010001110010",
						 "001001111111010001000100",
						 "001001111111010000010110",
						 "001001111111001111101000",
						 "001001111111001110111010",
						 "001001111111001110001100",
						 "001001111111001101011110",
						 "001001111111001100110000",
						 "001001111111001100000010",
						 "001001111111001011010100",
						 "001001111111001010100110",
						 "001001111111001001111000",
						 "001001111111001001001010",
						 "001001111111010011111100",
						 "001001111111010011001110",
						 "001001111111010010100000",
						 "001001111111010001110010",
						 "001001111111010001000100",
						 "001001111111010000010110",
						 "001001111111001111101000",
						 "001001111111001110111010",
						 "001001111111001110001100",
						 "001001111111001101011110",
						 "001001111111001100110000",
						 "001001111111001100000010",
						 "001001111111001011010100",
						 "001001111111001010100110",
						 "001001111111001001111000",
						 "001001111111001001001010",
						 "001001111111010100001011",
						 "001001111111010011011100",
						 "001001111111010010101101",
						 "001001111111010001111110",
						 "001001111111010001001111",
						 "001001111111010000100000",
						 "001001111111001111110001",
						 "001001111111001111000010",
						 "001001111111001110010011",
						 "001001111111001101100100",
						 "001001111111001100110101",
						 "001001111111001100000110",
						 "001001111111001011010111",
						 "001001111111001010101000",
						 "001001111111001001111001",
						 "001001111111001001001010",
						 "001001111111010100001011",
						 "001001111111010011011100",
						 "001001111111010010101101",
						 "001001111111010001111110",
						 "001001111111010001001111",
						 "001001111111010000100000",
						 "001001111111001111110001",
						 "001001111111001111000010",
						 "001001111111001110010011",
						 "001001111111001101100100",
						 "001001111111001100110101",
						 "001001111111001100000110",
						 "001001111111001011010111",
						 "001001111111001010101000",
						 "001001111111001001111001",
						 "001001111111001001001010",
						 "001001111100110001011100",
						 "001001111100110000101100",
						 "001001111100101111111100",
						 "001001111100101111001100",
						 "001001111100101110011100",
						 "001001111100101101101100",
						 "001001111100101100111100",
						 "001001111100101100001100",
						 "001001111100101011011100",
						 "001001111100101010101100",
						 "001001111100101001111100",
						 "001001111100101001001100",
						 "001001111100101000011100",
						 "001001111100100111101100",
						 "001001111100100110111100",
						 "001001111100100110001100",
						 "001001111100110001011100",
						 "001001111100110000101100",
						 "001001111100101111111100",
						 "001001111100101111001100",
						 "001001111100101110011100",
						 "001001111100101101101100",
						 "001001111100101100111100",
						 "001001111100101100001100",
						 "001001111100101011011100",
						 "001001111100101010101100",
						 "001001111100101001111100",
						 "001001111100101001001100",
						 "001001111100101000011100",
						 "001001111100100111101100",
						 "001001111100100110111100",
						 "001001111100100110001100",
						 "001001111100110001011100",
						 "001001111100110000101100",
						 "001001111100101111111100",
						 "001001111100101111001100",
						 "001001111100101110011100",
						 "001001111100101101101100",
						 "001001111100101100111100",
						 "001001111100101100001100",
						 "001001111100101011011100",
						 "001001111100101010101100",
						 "001001111100101001111100",
						 "001001111100101001001100",
						 "001001111100101000011100",
						 "001001111100100111101100",
						 "001001111100100110111100",
						 "001001111100100110001100",
						 "001001111100110001101011",
						 "001001111100110000111010",
						 "001001111100110000001001",
						 "001001111100101111011000",
						 "001001111100101110100111",
						 "001001111100101101110110",
						 "001001111100101101000101",
						 "001001111100101100010100",
						 "001001111100101011100011",
						 "001001111100101010110010",
						 "001001111100101010000001",
						 "001001111100101001010000",
						 "001001111100101000011111",
						 "001001111100100111101110",
						 "001001111100100110111101",
						 "001001111100100110001100",
						 "001001111100110001101011",
						 "001001111100110000111010",
						 "001001111100110000001001",
						 "001001111100101111011000",
						 "001001111100101110100111",
						 "001001111100101101110110",
						 "001001111100101101000101",
						 "001001111100101100010100",
						 "001001111100101011100011",
						 "001001111100101010110010",
						 "001001111100101010000001",
						 "001001111100101001010000",
						 "001001111100101000011111",
						 "001001111100100111101110",
						 "001001111100100110111101",
						 "001001111100100110001100",
						 "001001111100110001111010",
						 "001001111100110001001000",
						 "001001111100110000010110",
						 "001001111100101111100100",
						 "001001111100101110110010",
						 "001001111100101110000000",
						 "001001111100101101001110",
						 "001001111100101100011100",
						 "001001111100101011101010",
						 "001001111100101010111000",
						 "001001111100101010000110",
						 "001001111100101001010100",
						 "001001111100101000100010",
						 "001001111100100111110000",
						 "001001111100100110111110",
						 "001001111100100110001100",
						 "001001111100110001111010",
						 "001001111100110001001000",
						 "001001111100110000010110",
						 "001001111100101111100100",
						 "001001111100101110110010",
						 "001001111100101110000000",
						 "001001111100101101001110",
						 "001001111100101100011100",
						 "001001111100101011101010",
						 "001001111100101010111000",
						 "001001111100101010000110",
						 "001001111100101001010100",
						 "001001111100101000100010",
						 "001001111100100111110000",
						 "001001111100100110111110",
						 "001001111100100110001100",
						 "001001111100110001111010",
						 "001001111100110001001000",
						 "001001111100110000010110",
						 "001001111100101111100100",
						 "001001111100101110110010",
						 "001001111100101110000000",
						 "001001111100101101001110",
						 "001001111100101100011100",
						 "001001111100101011101010",
						 "001001111100101010111000",
						 "001001111100101010000110",
						 "001001111100101001010100",
						 "001001111100101000100010",
						 "001001111100100111110000",
						 "001001111100100110111110",
						 "001001111100100110001100",
						 "001001111100110010001001",
						 "001001111100110001010110",
						 "001001111100110000100011",
						 "001001111100101111110000",
						 "001001111100101110111101",
						 "001001111100101110001010",
						 "001001111100101101010111",
						 "001001111100101100100100",
						 "001001111100101011110001",
						 "001001111100101010111110",
						 "001001111100101010001011",
						 "001001111100101001011000",
						 "001001111100101000100101",
						 "001001111100100111110010",
						 "001001111100100110111111",
						 "001001111100100110001100",
						 "001001111100110010001001",
						 "001001111100110001010110",
						 "001001111100110000100011",
						 "001001111100101111110000",
						 "001001111100101110111101",
						 "001001111100101110001010",
						 "001001111100101101010111",
						 "001001111100101100100100",
						 "001001111100101011110001",
						 "001001111100101010111110",
						 "001001111100101010001011",
						 "001001111100101001011000",
						 "001001111100101000100101",
						 "001001111100100111110010",
						 "001001111100100110111111",
						 "001001111100100110001100",
						 "001001111100110010001001",
						 "001001111100110001010110",
						 "001001111100110000100011",
						 "001001111100101111110000",
						 "001001111100101110111101",
						 "001001111100101110001010",
						 "001001111100101101010111",
						 "001001111100101100100100",
						 "001001111100101011110001",
						 "001001111100101010111110",
						 "001001111100101010001011",
						 "001001111100101001011000",
						 "001001111100101000100101",
						 "001001111100100111110010",
						 "001001111100100110111111",
						 "001001111100100110001100",
						 "001001111100110010011000",
						 "001001111100110001100100",
						 "001001111100110000110000",
						 "001001111100101111111100",
						 "001001111100101111001000",
						 "001001111100101110010100",
						 "001001111100101101100000",
						 "001001111100101100101100",
						 "001001111100101011111000",
						 "001001111100101011000100",
						 "001001111100101010010000",
						 "001001111100101001011100",
						 "001001111100101000101000",
						 "001001111100100111110100",
						 "001001111100100111000000",
						 "001001111100100110001100",
						 "001001111100110010011000",
						 "001001111100110001100100",
						 "001001111100110000110000",
						 "001001111100101111111100",
						 "001001111100101111001000",
						 "001001111100101110010100",
						 "001001111100101101100000",
						 "001001111100101100101100",
						 "001001111100101011111000",
						 "001001111100101011000100",
						 "001001111100101010010000",
						 "001001111100101001011100",
						 "001001111100101000101000",
						 "001001111100100111110100",
						 "001001111100100111000000",
						 "001001111100100110001100",
						 "001001111010001111101001",
						 "001001111010001110110100",
						 "001001111010001101111111",
						 "001001111010001101001010",
						 "001001111010001100010101",
						 "001001111010001011100000",
						 "001001111010001010101011",
						 "001001111010001001110110",
						 "001001111010001001000001",
						 "001001111010001000001100",
						 "001001111010000111010111",
						 "001001111010000110100010",
						 "001001111010000101101101",
						 "001001111010000100111000",
						 "001001111010000100000011",
						 "001001111010000011001110",
						 "001001111010001111101001",
						 "001001111010001110110100",
						 "001001111010001101111111",
						 "001001111010001101001010",
						 "001001111010001100010101",
						 "001001111010001011100000",
						 "001001111010001010101011",
						 "001001111010001001110110",
						 "001001111010001001000001",
						 "001001111010001000001100",
						 "001001111010000111010111",
						 "001001111010000110100010",
						 "001001111010000101101101",
						 "001001111010000100111000",
						 "001001111010000100000011",
						 "001001111010000011001110",
						 "001001111010001111101001",
						 "001001111010001110110100",
						 "001001111010001101111111",
						 "001001111010001101001010",
						 "001001111010001100010101",
						 "001001111010001011100000",
						 "001001111010001010101011",
						 "001001111010001001110110",
						 "001001111010001001000001",
						 "001001111010001000001100",
						 "001001111010000111010111",
						 "001001111010000110100010",
						 "001001111010000101101101",
						 "001001111010000100111000",
						 "001001111010000100000011",
						 "001001111010000011001110",
						 "001001111010001111111000",
						 "001001111010001111000010",
						 "001001111010001110001100",
						 "001001111010001101010110",
						 "001001111010001100100000",
						 "001001111010001011101010",
						 "001001111010001010110100",
						 "001001111010001001111110",
						 "001001111010001001001000",
						 "001001111010001000010010",
						 "001001111010000111011100",
						 "001001111010000110100110",
						 "001001111010000101110000",
						 "001001111010000100111010",
						 "001001111010000100000100",
						 "001001111010000011001110",
						 "001001111010001111111000",
						 "001001111010001111000010",
						 "001001111010001110001100",
						 "001001111010001101010110",
						 "001001111010001100100000",
						 "001001111010001011101010",
						 "001001111010001010110100",
						 "001001111010001001111110",
						 "001001111010001001001000",
						 "001001111010001000010010",
						 "001001111010000111011100",
						 "001001111010000110100110",
						 "001001111010000101110000",
						 "001001111010000100111010",
						 "001001111010000100000100",
						 "001001111010000011001110",
						 "001001111010010000000111",
						 "001001111010001111010000",
						 "001001111010001110011001",
						 "001001111010001101100010",
						 "001001111010001100101011",
						 "001001111010001011110100",
						 "001001111010001010111101",
						 "001001111010001010000110",
						 "001001111010001001001111",
						 "001001111010001000011000",
						 "001001111010000111100001",
						 "001001111010000110101010",
						 "001001111010000101110011",
						 "001001111010000100111100",
						 "001001111010000100000101",
						 "001001111010000011001110",
						 "001001111010010000000111",
						 "001001111010001111010000",
						 "001001111010001110011001",
						 "001001111010001101100010",
						 "001001111010001100101011",
						 "001001111010001011110100",
						 "001001111010001010111101",
						 "001001111010001010000110",
						 "001001111010001001001111",
						 "001001111010001000011000",
						 "001001111010000111100001",
						 "001001111010000110101010",
						 "001001111010000101110011",
						 "001001111010000100111100",
						 "001001111010000100000101",
						 "001001111010000011001110",
						 "001001111010010000000111",
						 "001001111010001111010000",
						 "001001111010001110011001",
						 "001001111010001101100010",
						 "001001111010001100101011",
						 "001001111010001011110100",
						 "001001111010001010111101",
						 "001001111010001010000110",
						 "001001111010001001001111",
						 "001001111010001000011000",
						 "001001111010000111100001",
						 "001001111010000110101010",
						 "001001111010000101110011",
						 "001001111010000100111100",
						 "001001111010000100000101",
						 "001001111010000011001110",
						 "001001111010010000010110",
						 "001001111010001111011110",
						 "001001111010001110100110",
						 "001001111010001101101110",
						 "001001111010001100110110",
						 "001001111010001011111110",
						 "001001111010001011000110",
						 "001001111010001010001110",
						 "001001111010001001010110",
						 "001001111010001000011110",
						 "001001111010000111100110",
						 "001001111010000110101110",
						 "001001111010000101110110",
						 "001001111010000100111110",
						 "001001111010000100000110",
						 "001001111010000011001110",
						 "001001111010010000010110",
						 "001001111010001111011110",
						 "001001111010001110100110",
						 "001001111010001101101110",
						 "001001111010001100110110",
						 "001001111010001011111110",
						 "001001111010001011000110",
						 "001001111010001010001110",
						 "001001111010001001010110",
						 "001001111010001000011110",
						 "001001111010000111100110",
						 "001001111010000110101110",
						 "001001111010000101110110",
						 "001001111010000100111110",
						 "001001111010000100000110",
						 "001001111010000011001110",
						 "001001111010010000010110",
						 "001001111010001111011110",
						 "001001111010001110100110",
						 "001001111010001101101110",
						 "001001111010001100110110",
						 "001001111010001011111110",
						 "001001111010001011000110",
						 "001001111010001010001110",
						 "001001111010001001010110",
						 "001001111010001000011110",
						 "001001111010000111100110",
						 "001001111010000110101110",
						 "001001111010000101110110",
						 "001001111010000100111110",
						 "001001111010000100000110",
						 "001001111010000011001110",
						 "001001111010010000100101",
						 "001001111010001111101100",
						 "001001111010001110110011",
						 "001001111010001101111010",
						 "001001111010001101000001",
						 "001001111010001100001000",
						 "001001111010001011001111",
						 "001001111010001010010110",
						 "001001111010001001011101",
						 "001001111010001000100100",
						 "001001111010000111101011",
						 "001001111010000110110010",
						 "001001111010000101111001",
						 "001001111010000101000000",
						 "001001111010000100000111",
						 "001001111010000011001110",
						 "001001110111101101100111",
						 "001001110111101100101110",
						 "001001110111101011110101",
						 "001001110111101010111100",
						 "001001110111101010000011",
						 "001001110111101001001010",
						 "001001110111101000010001",
						 "001001110111100111011000",
						 "001001110111100110011111",
						 "001001110111100101100110",
						 "001001110111100100101101",
						 "001001110111100011110100",
						 "001001110111100010111011",
						 "001001110111100010000010",
						 "001001110111100001001001",
						 "001001110111100000010000",
						 "001001110111101101110110",
						 "001001110111101100111100",
						 "001001110111101100000010",
						 "001001110111101011001000",
						 "001001110111101010001110",
						 "001001110111101001010100",
						 "001001110111101000011010",
						 "001001110111100111100000",
						 "001001110111100110100110",
						 "001001110111100101101100",
						 "001001110111100100110010",
						 "001001110111100011111000",
						 "001001110111100010111110",
						 "001001110111100010000100",
						 "001001110111100001001010",
						 "001001110111100000010000",
						 "001001110111101101110110",
						 "001001110111101100111100",
						 "001001110111101100000010",
						 "001001110111101011001000",
						 "001001110111101010001110",
						 "001001110111101001010100",
						 "001001110111101000011010",
						 "001001110111100111100000",
						 "001001110111100110100110",
						 "001001110111100101101100",
						 "001001110111100100110010",
						 "001001110111100011111000",
						 "001001110111100010111110",
						 "001001110111100010000100",
						 "001001110111100001001010",
						 "001001110111100000010000",
						 "001001110111101101110110",
						 "001001110111101100111100",
						 "001001110111101100000010",
						 "001001110111101011001000",
						 "001001110111101010001110",
						 "001001110111101001010100",
						 "001001110111101000011010",
						 "001001110111100111100000",
						 "001001110111100110100110",
						 "001001110111100101101100",
						 "001001110111100100110010",
						 "001001110111100011111000",
						 "001001110111100010111110",
						 "001001110111100010000100",
						 "001001110111100001001010",
						 "001001110111100000010000",
						 "001001110111101110000101",
						 "001001110111101101001010",
						 "001001110111101100001111",
						 "001001110111101011010100",
						 "001001110111101010011001",
						 "001001110111101001011110",
						 "001001110111101000100011",
						 "001001110111100111101000",
						 "001001110111100110101101",
						 "001001110111100101110010",
						 "001001110111100100110111",
						 "001001110111100011111100",
						 "001001110111100011000001",
						 "001001110111100010000110",
						 "001001110111100001001011",
						 "001001110111100000010000",
						 "001001110111101110000101",
						 "001001110111101101001010",
						 "001001110111101100001111",
						 "001001110111101011010100",
						 "001001110111101010011001",
						 "001001110111101001011110",
						 "001001110111101000100011",
						 "001001110111100111101000",
						 "001001110111100110101101",
						 "001001110111100101110010",
						 "001001110111100100110111",
						 "001001110111100011111100",
						 "001001110111100011000001",
						 "001001110111100010000110",
						 "001001110111100001001011",
						 "001001110111100000010000",
						 "001001110111101110000101",
						 "001001110111101101001010",
						 "001001110111101100001111",
						 "001001110111101011010100",
						 "001001110111101010011001",
						 "001001110111101001011110",
						 "001001110111101000100011",
						 "001001110111100111101000",
						 "001001110111100110101101",
						 "001001110111100101110010",
						 "001001110111100100110111",
						 "001001110111100011111100",
						 "001001110111100011000001",
						 "001001110111100010000110",
						 "001001110111100001001011",
						 "001001110111100000010000",
						 "001001110111101110010100",
						 "001001110111101101011000",
						 "001001110111101100011100",
						 "001001110111101011100000",
						 "001001110111101010100100",
						 "001001110111101001101000",
						 "001001110111101000101100",
						 "001001110111100111110000",
						 "001001110111100110110100",
						 "001001110111100101111000",
						 "001001110111100100111100",
						 "001001110111100100000000",
						 "001001110111100011000100",
						 "001001110111100010001000",
						 "001001110111100001001100",
						 "001001110111100000010000",
						 "001001110111101110010100",
						 "001001110111101101011000",
						 "001001110111101100011100",
						 "001001110111101011100000",
						 "001001110111101010100100",
						 "001001110111101001101000",
						 "001001110111101000101100",
						 "001001110111100111110000",
						 "001001110111100110110100",
						 "001001110111100101111000",
						 "001001110111100100111100",
						 "001001110111100100000000",
						 "001001110111100011000100",
						 "001001110111100010001000",
						 "001001110111100001001100",
						 "001001110111100000010000",
						 "001001110111101110100011",
						 "001001110111101101100110",
						 "001001110111101100101001",
						 "001001110111101011101100",
						 "001001110111101010101111",
						 "001001110111101001110010",
						 "001001110111101000110101",
						 "001001110111100111111000",
						 "001001110111100110111011",
						 "001001110111100101111110",
						 "001001110111100101000001",
						 "001001110111100100000100",
						 "001001110111100011000111",
						 "001001110111100010001010",
						 "001001110111100001001101",
						 "001001110111100000010000",
						 "001001110111101110100011",
						 "001001110111101101100110",
						 "001001110111101100101001",
						 "001001110111101011101100",
						 "001001110111101010101111",
						 "001001110111101001110010",
						 "001001110111101000110101",
						 "001001110111100111111000",
						 "001001110111100110111011",
						 "001001110111100101111110",
						 "001001110111100101000001",
						 "001001110111100100000100",
						 "001001110111100011000111",
						 "001001110111100010001010",
						 "001001110111100001001101",
						 "001001110111100000010000",
						 "001001110101001011100101",
						 "001001110101001010101000",
						 "001001110101001001101011",
						 "001001110101001000101110",
						 "001001110101000111110001",
						 "001001110101000110110100",
						 "001001110101000101110111",
						 "001001110101000100111010",
						 "001001110101000011111101",
						 "001001110101000011000000",
						 "001001110101000010000011",
						 "001001110101000001000110",
						 "001001110101000000001001",
						 "001001110100111111001100",
						 "001001110100111110001111",
						 "001001110100111101010010",
						 "001001110101001011110100",
						 "001001110101001010110110",
						 "001001110101001001111000",
						 "001001110101001000111010",
						 "001001110101000111111100",
						 "001001110101000110111110",
						 "001001110101000110000000",
						 "001001110101000101000010",
						 "001001110101000100000100",
						 "001001110101000011000110",
						 "001001110101000010001000",
						 "001001110101000001001010",
						 "001001110101000000001100",
						 "001001110100111111001110",
						 "001001110100111110010000",
						 "001001110100111101010010",
						 "001001110101001011110100",
						 "001001110101001010110110",
						 "001001110101001001111000",
						 "001001110101001000111010",
						 "001001110101000111111100",
						 "001001110101000110111110",
						 "001001110101000110000000",
						 "001001110101000101000010",
						 "001001110101000100000100",
						 "001001110101000011000110",
						 "001001110101000010001000",
						 "001001110101000001001010",
						 "001001110101000000001100",
						 "001001110100111111001110",
						 "001001110100111110010000",
						 "001001110100111101010010",
						 "001001110101001100000011",
						 "001001110101001011000100",
						 "001001110101001010000101",
						 "001001110101001001000110",
						 "001001110101001000000111",
						 "001001110101000111001000",
						 "001001110101000110001001",
						 "001001110101000101001010",
						 "001001110101000100001011",
						 "001001110101000011001100",
						 "001001110101000010001101",
						 "001001110101000001001110",
						 "001001110101000000001111",
						 "001001110100111111010000",
						 "001001110100111110010001",
						 "001001110100111101010010",
						 "001001110101001100000011",
						 "001001110101001011000100",
						 "001001110101001010000101",
						 "001001110101001001000110",
						 "001001110101001000000111",
						 "001001110101000111001000",
						 "001001110101000110001001",
						 "001001110101000101001010",
						 "001001110101000100001011",
						 "001001110101000011001100",
						 "001001110101000010001101",
						 "001001110101000001001110",
						 "001001110101000000001111",
						 "001001110100111111010000",
						 "001001110100111110010001",
						 "001001110100111101010010",
						 "001001110101001100000011",
						 "001001110101001011000100",
						 "001001110101001010000101",
						 "001001110101001001000110",
						 "001001110101001000000111",
						 "001001110101000111001000",
						 "001001110101000110001001",
						 "001001110101000101001010",
						 "001001110101000100001011",
						 "001001110101000011001100",
						 "001001110101000010001101",
						 "001001110101000001001110",
						 "001001110101000000001111",
						 "001001110100111111010000",
						 "001001110100111110010001",
						 "001001110100111101010010",
						 "001001110101001100010010",
						 "001001110101001011010010",
						 "001001110101001010010010",
						 "001001110101001001010010",
						 "001001110101001000010010",
						 "001001110101000111010010",
						 "001001110101000110010010",
						 "001001110101000101010010",
						 "001001110101000100010010",
						 "001001110101000011010010",
						 "001001110101000010010010",
						 "001001110101000001010010",
						 "001001110101000000010010",
						 "001001110100111111010010",
						 "001001110100111110010010",
						 "001001110100111101010010",
						 "001001110101001100010010",
						 "001001110101001011010010",
						 "001001110101001010010010",
						 "001001110101001001010010",
						 "001001110101001000010010",
						 "001001110101000111010010",
						 "001001110101000110010010",
						 "001001110101000101010010",
						 "001001110101000100010010",
						 "001001110101000011010010",
						 "001001110101000010010010",
						 "001001110101000001010010",
						 "001001110101000000010010",
						 "001001110100111111010010",
						 "001001110100111110010010",
						 "001001110100111101010010",
						 "001001110101001100010010",
						 "001001110101001011010010",
						 "001001110101001010010010",
						 "001001110101001001010010",
						 "001001110101001000010010",
						 "001001110101000111010010",
						 "001001110101000110010010",
						 "001001110101000101010010",
						 "001001110101000100010010",
						 "001001110101000011010010",
						 "001001110101000010010010",
						 "001001110101000001010010",
						 "001001110101000000010010",
						 "001001110100111111010010",
						 "001001110100111110010010",
						 "001001110100111101010010",
						 "001001110101001100100001",
						 "001001110101001011100000",
						 "001001110101001010011111",
						 "001001110101001001011110",
						 "001001110101001000011101",
						 "001001110101000111011100",
						 "001001110101000110011011",
						 "001001110101000101011010",
						 "001001110101000100011001",
						 "001001110101000011011000",
						 "001001110101000010010111",
						 "001001110101000001010110",
						 "001001110101000000010101",
						 "001001110100111111010100",
						 "001001110100111110010011",
						 "001001110100111101010010",
						 "001001110010101001100011",
						 "001001110010101000100010",
						 "001001110010100111100001",
						 "001001110010100110100000",
						 "001001110010100101011111",
						 "001001110010100100011110",
						 "001001110010100011011101",
						 "001001110010100010011100",
						 "001001110010100001011011",
						 "001001110010100000011010",
						 "001001110010011111011001",
						 "001001110010011110011000",
						 "001001110010011101010111",
						 "001001110010011100010110",
						 "001001110010011011010101",
						 "001001110010011010010100",
						 "001001110010101001110010",
						 "001001110010101000110000",
						 "001001110010100111101110",
						 "001001110010100110101100",
						 "001001110010100101101010",
						 "001001110010100100101000",
						 "001001110010100011100110",
						 "001001110010100010100100",
						 "001001110010100001100010",
						 "001001110010100000100000",
						 "001001110010011111011110",
						 "001001110010011110011100",
						 "001001110010011101011010",
						 "001001110010011100011000",
						 "001001110010011011010110",
						 "001001110010011010010100",
						 "001001110010101001110010",
						 "001001110010101000110000",
						 "001001110010100111101110",
						 "001001110010100110101100",
						 "001001110010100101101010",
						 "001001110010100100101000",
						 "001001110010100011100110",
						 "001001110010100010100100",
						 "001001110010100001100010",
						 "001001110010100000100000",
						 "001001110010011111011110",
						 "001001110010011110011100",
						 "001001110010011101011010",
						 "001001110010011100011000",
						 "001001110010011011010110",
						 "001001110010011010010100",
						 "001001110010101001110010",
						 "001001110010101000110000",
						 "001001110010100111101110",
						 "001001110010100110101100",
						 "001001110010100101101010",
						 "001001110010100100101000",
						 "001001110010100011100110",
						 "001001110010100010100100",
						 "001001110010100001100010",
						 "001001110010100000100000",
						 "001001110010011111011110",
						 "001001110010011110011100",
						 "001001110010011101011010",
						 "001001110010011100011000",
						 "001001110010011011010110",
						 "001001110010011010010100",
						 "001001110010101010000001",
						 "001001110010101000111110",
						 "001001110010100111111011",
						 "001001110010100110111000",
						 "001001110010100101110101",
						 "001001110010100100110010",
						 "001001110010100011101111",
						 "001001110010100010101100",
						 "001001110010100001101001",
						 "001001110010100000100110",
						 "001001110010011111100011",
						 "001001110010011110100000",
						 "001001110010011101011101",
						 "001001110010011100011010",
						 "001001110010011011010111",
						 "001001110010011010010100",
						 "001001110010101010000001",
						 "001001110010101000111110",
						 "001001110010100111111011",
						 "001001110010100110111000",
						 "001001110010100101110101",
						 "001001110010100100110010",
						 "001001110010100011101111",
						 "001001110010100010101100",
						 "001001110010100001101001",
						 "001001110010100000100110",
						 "001001110010011111100011",
						 "001001110010011110100000",
						 "001001110010011101011101",
						 "001001110010011100011010",
						 "001001110010011011010111",
						 "001001110010011010010100",
						 "001001110010101010000001",
						 "001001110010101000111110",
						 "001001110010100111111011",
						 "001001110010100110111000",
						 "001001110010100101110101",
						 "001001110010100100110010",
						 "001001110010100011101111",
						 "001001110010100010101100",
						 "001001110010100001101001",
						 "001001110010100000100110",
						 "001001110010011111100011",
						 "001001110010011110100000",
						 "001001110010011101011101",
						 "001001110010011100011010",
						 "001001110010011011010111",
						 "001001110010011010010100",
						 "001001110010101010010000",
						 "001001110010101001001100",
						 "001001110010101000001000",
						 "001001110010100111000100",
						 "001001110010100110000000",
						 "001001110010100100111100",
						 "001001110010100011111000",
						 "001001110010100010110100",
						 "001001110010100001110000",
						 "001001110010100000101100",
						 "001001110010011111101000",
						 "001001110010011110100100",
						 "001001110010011101100000",
						 "001001110010011100011100",
						 "001001110010011011011000",
						 "001001110010011010010100",
						 "001001110010101010010000",
						 "001001110010101001001100",
						 "001001110010101000001000",
						 "001001110010100111000100",
						 "001001110010100110000000",
						 "001001110010100100111100",
						 "001001110010100011111000",
						 "001001110010100010110100",
						 "001001110010100001110000",
						 "001001110010100000101100",
						 "001001110010011111101000",
						 "001001110010011110100100",
						 "001001110010011101100000",
						 "001001110010011100011100",
						 "001001110010011011011000",
						 "001001110010011010010100",
						 "001001110010101010011111",
						 "001001110010101001011010",
						 "001001110010101000010101",
						 "001001110010100111010000",
						 "001001110010100110001011",
						 "001001110010100101000110",
						 "001001110010100100000001",
						 "001001110010100010111100",
						 "001001110010100001110111",
						 "001001110010100000110010",
						 "001001110010011111101101",
						 "001001110010011110101000",
						 "001001110010011101100011",
						 "001001110010011100011110",
						 "001001110010011011011001",
						 "001001110010011010010100",
						 "001001110000000111100001",
						 "001001110000000110011100",
						 "001001110000000101010111",
						 "001001110000000100010010",
						 "001001110000000011001101",
						 "001001110000000010001000",
						 "001001110000000001000011",
						 "001001101111111111111110",
						 "001001101111111110111001",
						 "001001101111111101110100",
						 "001001101111111100101111",
						 "001001101111111011101010",
						 "001001101111111010100101",
						 "001001101111111001100000",
						 "001001101111111000011011",
						 "001001101111110111010110",
						 "001001110000000111100001",
						 "001001110000000110011100",
						 "001001110000000101010111",
						 "001001110000000100010010",
						 "001001110000000011001101",
						 "001001110000000010001000",
						 "001001110000000001000011",
						 "001001101111111111111110",
						 "001001101111111110111001",
						 "001001101111111101110100",
						 "001001101111111100101111",
						 "001001101111111011101010",
						 "001001101111111010100101",
						 "001001101111111001100000",
						 "001001101111111000011011",
						 "001001101111110111010110",
						 "001001110000000111110000",
						 "001001110000000110101010",
						 "001001110000000101100100",
						 "001001110000000100011110",
						 "001001110000000011011000",
						 "001001110000000010010010",
						 "001001110000000001001100",
						 "001001110000000000000110",
						 "001001101111111111000000",
						 "001001101111111101111010",
						 "001001101111111100110100",
						 "001001101111111011101110",
						 "001001101111111010101000",
						 "001001101111111001100010",
						 "001001101111111000011100",
						 "001001101111110111010110",
						 "001001110000000111110000",
						 "001001110000000110101010",
						 "001001110000000101100100",
						 "001001110000000100011110",
						 "001001110000000011011000",
						 "001001110000000010010010",
						 "001001110000000001001100",
						 "001001110000000000000110",
						 "001001101111111111000000",
						 "001001101111111101111010",
						 "001001101111111100110100",
						 "001001101111111011101110",
						 "001001101111111010101000",
						 "001001101111111001100010",
						 "001001101111111000011100",
						 "001001101111110111010110",
						 "001001110000000111110000",
						 "001001110000000110101010",
						 "001001110000000101100100",
						 "001001110000000100011110",
						 "001001110000000011011000",
						 "001001110000000010010010",
						 "001001110000000001001100",
						 "001001110000000000000110",
						 "001001101111111111000000",
						 "001001101111111101111010",
						 "001001101111111100110100",
						 "001001101111111011101110",
						 "001001101111111010101000",
						 "001001101111111001100010",
						 "001001101111111000011100",
						 "001001101111110111010110",
						 "001001110000000111111111",
						 "001001110000000110111000",
						 "001001110000000101110001",
						 "001001110000000100101010",
						 "001001110000000011100011",
						 "001001110000000010011100",
						 "001001110000000001010101",
						 "001001110000000000001110",
						 "001001101111111111000111",
						 "001001101111111110000000",
						 "001001101111111100111001",
						 "001001101111111011110010",
						 "001001101111111010101011",
						 "001001101111111001100100",
						 "001001101111111000011101",
						 "001001101111110111010110",
						 "001001110000000111111111",
						 "001001110000000110111000",
						 "001001110000000101110001",
						 "001001110000000100101010",
						 "001001110000000011100011",
						 "001001110000000010011100",
						 "001001110000000001010101",
						 "001001110000000000001110",
						 "001001101111111111000111",
						 "001001101111111110000000",
						 "001001101111111100111001",
						 "001001101111111011110010",
						 "001001101111111010101011",
						 "001001101111111001100100",
						 "001001101111111000011101",
						 "001001101111110111010110",
						 "001001110000001000001110",
						 "001001110000000111000110",
						 "001001110000000101111110",
						 "001001110000000100110110",
						 "001001110000000011101110",
						 "001001110000000010100110",
						 "001001110000000001011110",
						 "001001110000000000010110",
						 "001001101111111111001110",
						 "001001101111111110000110",
						 "001001101111111100111110",
						 "001001101111111011110110",
						 "001001101111111010101110",
						 "001001101111111001100110",
						 "001001101111111000011110",
						 "001001101111110111010110",
						 "001001110000001000001110",
						 "001001110000000111000110",
						 "001001110000000101111110",
						 "001001110000000100110110",
						 "001001110000000011101110",
						 "001001110000000010100110",
						 "001001110000000001011110",
						 "001001110000000000010110",
						 "001001101111111111001110",
						 "001001101111111110000110",
						 "001001101111111100111110",
						 "001001101111111011110110",
						 "001001101111111010101110",
						 "001001101111111001100110",
						 "001001101111111000011110",
						 "001001101111110111010110",
						 "001001101101100101010000",
						 "001001101101100100001000",
						 "001001101101100011000000",
						 "001001101101100001111000",
						 "001001101101100000110000",
						 "001001101101011111101000",
						 "001001101101011110100000",
						 "001001101101011101011000",
						 "001001101101011100010000",
						 "001001101101011011001000",
						 "001001101101011010000000",
						 "001001101101011000111000",
						 "001001101101010111110000",
						 "001001101101010110101000",
						 "001001101101010101100000",
						 "001001101101010100011000",
						 "001001101101100101011111",
						 "001001101101100100010110",
						 "001001101101100011001101",
						 "001001101101100010000100",
						 "001001101101100000111011",
						 "001001101101011111110010",
						 "001001101101011110101001",
						 "001001101101011101100000",
						 "001001101101011100010111",
						 "001001101101011011001110",
						 "001001101101011010000101",
						 "001001101101011000111100",
						 "001001101101010111110011",
						 "001001101101010110101010",
						 "001001101101010101100001",
						 "001001101101010100011000",
						 "001001101101100101011111",
						 "001001101101100100010110",
						 "001001101101100011001101",
						 "001001101101100010000100",
						 "001001101101100000111011",
						 "001001101101011111110010",
						 "001001101101011110101001",
						 "001001101101011101100000",
						 "001001101101011100010111",
						 "001001101101011011001110",
						 "001001101101011010000101",
						 "001001101101011000111100",
						 "001001101101010111110011",
						 "001001101101010110101010",
						 "001001101101010101100001",
						 "001001101101010100011000",
						 "001001101101100101011111",
						 "001001101101100100010110",
						 "001001101101100011001101",
						 "001001101101100010000100",
						 "001001101101100000111011",
						 "001001101101011111110010",
						 "001001101101011110101001",
						 "001001101101011101100000",
						 "001001101101011100010111",
						 "001001101101011011001110",
						 "001001101101011010000101",
						 "001001101101011000111100",
						 "001001101101010111110011",
						 "001001101101010110101010",
						 "001001101101010101100001",
						 "001001101101010100011000",
						 "001001101101100101101110",
						 "001001101101100100100100",
						 "001001101101100011011010",
						 "001001101101100010010000",
						 "001001101101100001000110",
						 "001001101101011111111100",
						 "001001101101011110110010",
						 "001001101101011101101000",
						 "001001101101011100011110",
						 "001001101101011011010100",
						 "001001101101011010001010",
						 "001001101101011001000000",
						 "001001101101010111110110",
						 "001001101101010110101100",
						 "001001101101010101100010",
						 "001001101101010100011000",
						 "001001101101100101101110",
						 "001001101101100100100100",
						 "001001101101100011011010",
						 "001001101101100010010000",
						 "001001101101100001000110",
						 "001001101101011111111100",
						 "001001101101011110110010",
						 "001001101101011101101000",
						 "001001101101011100011110",
						 "001001101101011011010100",
						 "001001101101011010001010",
						 "001001101101011001000000",
						 "001001101101010111110110",
						 "001001101101010110101100",
						 "001001101101010101100010",
						 "001001101101010100011000",
						 "001001101101100101111101",
						 "001001101101100100110010",
						 "001001101101100011100111",
						 "001001101101100010011100",
						 "001001101101100001010001",
						 "001001101101100000000110",
						 "001001101101011110111011",
						 "001001101101011101110000",
						 "001001101101011100100101",
						 "001001101101011011011010",
						 "001001101101011010001111",
						 "001001101101011001000100",
						 "001001101101010111111001",
						 "001001101101010110101110",
						 "001001101101010101100011",
						 "001001101101010100011000",
						 "001001101101100101111101",
						 "001001101101100100110010",
						 "001001101101100011100111",
						 "001001101101100010011100",
						 "001001101101100001010001",
						 "001001101101100000000110",
						 "001001101101011110111011",
						 "001001101101011101110000",
						 "001001101101011100100101",
						 "001001101101011011011010",
						 "001001101101011010001111",
						 "001001101101011001000100",
						 "001001101101010111111001",
						 "001001101101010110101110",
						 "001001101101010101100011",
						 "001001101101010100011000",
						 "001001101101100101111101",
						 "001001101101100100110010",
						 "001001101101100011100111",
						 "001001101101100010011100",
						 "001001101101100001010001",
						 "001001101101100000000110",
						 "001001101101011110111011",
						 "001001101101011101110000",
						 "001001101101011100100101",
						 "001001101101011011011010",
						 "001001101101011010001111",
						 "001001101101011001000100",
						 "001001101101010111111001",
						 "001001101101010110101110",
						 "001001101101010101100011",
						 "001001101101010100011000",
						 "001001101011000011001110",
						 "001001101011000010000010",
						 "001001101011000000110110",
						 "001001101010111111101010",
						 "001001101010111110011110",
						 "001001101010111101010010",
						 "001001101010111100000110",
						 "001001101010111010111010",
						 "001001101010111001101110",
						 "001001101010111000100010",
						 "001001101010110111010110",
						 "001001101010110110001010",
						 "001001101010110100111110",
						 "001001101010110011110010",
						 "001001101010110010100110",
						 "001001101010110001011010",
						 "001001101011000011001110",
						 "001001101011000010000010",
						 "001001101011000000110110",
						 "001001101010111111101010",
						 "001001101010111110011110",
						 "001001101010111101010010",
						 "001001101010111100000110",
						 "001001101010111010111010",
						 "001001101010111001101110",
						 "001001101010111000100010",
						 "001001101010110111010110",
						 "001001101010110110001010",
						 "001001101010110100111110",
						 "001001101010110011110010",
						 "001001101010110010100110",
						 "001001101010110001011010",
						 "001001101011000011001110",
						 "001001101011000010000010",
						 "001001101011000000110110",
						 "001001101010111111101010",
						 "001001101010111110011110",
						 "001001101010111101010010",
						 "001001101010111100000110",
						 "001001101010111010111010",
						 "001001101010111001101110",
						 "001001101010111000100010",
						 "001001101010110111010110",
						 "001001101010110110001010",
						 "001001101010110100111110",
						 "001001101010110011110010",
						 "001001101010110010100110",
						 "001001101010110001011010",
						 "001001101011000011011101",
						 "001001101011000010010000",
						 "001001101011000001000011",
						 "001001101010111111110110",
						 "001001101010111110101001",
						 "001001101010111101011100",
						 "001001101010111100001111",
						 "001001101010111011000010",
						 "001001101010111001110101",
						 "001001101010111000101000",
						 "001001101010110111011011",
						 "001001101010110110001110",
						 "001001101010110101000001",
						 "001001101010110011110100",
						 "001001101010110010100111",
						 "001001101010110001011010",
						 "001001101011000011011101",
						 "001001101011000010010000",
						 "001001101011000001000011",
						 "001001101010111111110110",
						 "001001101010111110101001",
						 "001001101010111101011100",
						 "001001101010111100001111",
						 "001001101010111011000010",
						 "001001101010111001110101",
						 "001001101010111000101000",
						 "001001101010110111011011",
						 "001001101010110110001110",
						 "001001101010110101000001",
						 "001001101010110011110100",
						 "001001101010110010100111",
						 "001001101010110001011010",
						 "001001101011000011101100",
						 "001001101011000010011110",
						 "001001101011000001010000",
						 "001001101011000000000010",
						 "001001101010111110110100",
						 "001001101010111101100110",
						 "001001101010111100011000",
						 "001001101010111011001010",
						 "001001101010111001111100",
						 "001001101010111000101110",
						 "001001101010110111100000",
						 "001001101010110110010010",
						 "001001101010110101000100",
						 "001001101010110011110110",
						 "001001101010110010101000",
						 "001001101010110001011010",
						 "001001101011000011101100",
						 "001001101011000010011110",
						 "001001101011000001010000",
						 "001001101011000000000010",
						 "001001101010111110110100",
						 "001001101010111101100110",
						 "001001101010111100011000",
						 "001001101010111011001010",
						 "001001101010111001111100",
						 "001001101010111000101110",
						 "001001101010110111100000",
						 "001001101010110110010010",
						 "001001101010110101000100",
						 "001001101010110011110110",
						 "001001101010110010101000",
						 "001001101010110001011010",
						 "001001101011000011101100",
						 "001001101011000010011110",
						 "001001101011000001010000",
						 "001001101011000000000010",
						 "001001101010111110110100",
						 "001001101010111101100110",
						 "001001101010111100011000",
						 "001001101010111011001010",
						 "001001101010111001111100",
						 "001001101010111000101110",
						 "001001101010110111100000",
						 "001001101010110110010010",
						 "001001101010110101000100",
						 "001001101010110011110110",
						 "001001101010110010101000",
						 "001001101010110001011010",
						 "001001101000100000111101",
						 "001001101000011111101110",
						 "001001101000011110011111",
						 "001001101000011101010000",
						 "001001101000011100000001",
						 "001001101000011010110010",
						 "001001101000011001100011",
						 "001001101000011000010100",
						 "001001101000010111000101",
						 "001001101000010101110110",
						 "001001101000010100100111",
						 "001001101000010011011000",
						 "001001101000010010001001",
						 "001001101000010000111010",
						 "001001101000001111101011",
						 "001001101000001110011100",
						 "001001101000100000111101",
						 "001001101000011111101110",
						 "001001101000011110011111",
						 "001001101000011101010000",
						 "001001101000011100000001",
						 "001001101000011010110010",
						 "001001101000011001100011",
						 "001001101000011000010100",
						 "001001101000010111000101",
						 "001001101000010101110110",
						 "001001101000010100100111",
						 "001001101000010011011000",
						 "001001101000010010001001",
						 "001001101000010000111010",
						 "001001101000001111101011",
						 "001001101000001110011100",
						 "001001101000100000111101",
						 "001001101000011111101110",
						 "001001101000011110011111",
						 "001001101000011101010000",
						 "001001101000011100000001",
						 "001001101000011010110010",
						 "001001101000011001100011",
						 "001001101000011000010100",
						 "001001101000010111000101",
						 "001001101000010101110110",
						 "001001101000010100100111",
						 "001001101000010011011000",
						 "001001101000010010001001",
						 "001001101000010000111010",
						 "001001101000001111101011",
						 "001001101000001110011100",
						 "001001101000100001001100",
						 "001001101000011111111100",
						 "001001101000011110101100",
						 "001001101000011101011100",
						 "001001101000011100001100",
						 "001001101000011010111100",
						 "001001101000011001101100",
						 "001001101000011000011100",
						 "001001101000010111001100",
						 "001001101000010101111100",
						 "001001101000010100101100",
						 "001001101000010011011100",
						 "001001101000010010001100",
						 "001001101000010000111100",
						 "001001101000001111101100",
						 "001001101000001110011100",
						 "001001101000100001001100",
						 "001001101000011111111100",
						 "001001101000011110101100",
						 "001001101000011101011100",
						 "001001101000011100001100",
						 "001001101000011010111100",
						 "001001101000011001101100",
						 "001001101000011000011100",
						 "001001101000010111001100",
						 "001001101000010101111100",
						 "001001101000010100101100",
						 "001001101000010011011100",
						 "001001101000010010001100",
						 "001001101000010000111100",
						 "001001101000001111101100",
						 "001001101000001110011100",
						 "001001101000100001011011",
						 "001001101000100000001010",
						 "001001101000011110111001",
						 "001001101000011101101000",
						 "001001101000011100010111",
						 "001001101000011011000110",
						 "001001101000011001110101",
						 "001001101000011000100100",
						 "001001101000010111010011",
						 "001001101000010110000010",
						 "001001101000010100110001",
						 "001001101000010011100000",
						 "001001101000010010001111",
						 "001001101000010000111110",
						 "001001101000001111101101",
						 "001001101000001110011100",
						 "001001101000100001011011",
						 "001001101000100000001010",
						 "001001101000011110111001",
						 "001001101000011101101000",
						 "001001101000011100010111",
						 "001001101000011011000110",
						 "001001101000011001110101",
						 "001001101000011000100100",
						 "001001101000010111010011",
						 "001001101000010110000010",
						 "001001101000010100110001",
						 "001001101000010011100000",
						 "001001101000010010001111",
						 "001001101000010000111110",
						 "001001101000001111101101",
						 "001001101000001110011100",
						 "001001101000100001011011",
						 "001001101000100000001010",
						 "001001101000011110111001",
						 "001001101000011101101000",
						 "001001101000011100010111",
						 "001001101000011011000110",
						 "001001101000011001110101",
						 "001001101000011000100100",
						 "001001101000010111010011",
						 "001001101000010110000010",
						 "001001101000010100110001",
						 "001001101000010011100000",
						 "001001101000010010001111",
						 "001001101000010000111110",
						 "001001101000001111101101",
						 "001001101000001110011100",
						 "001001101000100001101010",
						 "001001101000100000011000",
						 "001001101000011111000110",
						 "001001101000011101110100",
						 "001001101000011100100010",
						 "001001101000011011010000",
						 "001001101000011001111110",
						 "001001101000011000101100",
						 "001001101000010111011010",
						 "001001101000010110001000",
						 "001001101000010100110110",
						 "001001101000010011100100",
						 "001001101000010010010010",
						 "001001101000010001000000",
						 "001001101000001111101110",
						 "001001101000001110011100",
						 "001001100101111110101100",
						 "001001100101111101011010",
						 "001001100101111100001000",
						 "001001100101111010110110",
						 "001001100101111001100100",
						 "001001100101111000010010",
						 "001001100101110111000000",
						 "001001100101110101101110",
						 "001001100101110100011100",
						 "001001100101110011001010",
						 "001001100101110001111000",
						 "001001100101110000100110",
						 "001001100101101111010100",
						 "001001100101101110000010",
						 "001001100101101100110000",
						 "001001100101101011011110",
						 "001001100101111110101100",
						 "001001100101111101011010",
						 "001001100101111100001000",
						 "001001100101111010110110",
						 "001001100101111001100100",
						 "001001100101111000010010",
						 "001001100101110111000000",
						 "001001100101110101101110",
						 "001001100101110100011100",
						 "001001100101110011001010",
						 "001001100101110001111000",
						 "001001100101110000100110",
						 "001001100101101111010100",
						 "001001100101101110000010",
						 "001001100101101100110000",
						 "001001100101101011011110",
						 "001001100101111110111011",
						 "001001100101111101101000",
						 "001001100101111100010101",
						 "001001100101111011000010",
						 "001001100101111001101111",
						 "001001100101111000011100",
						 "001001100101110111001001",
						 "001001100101110101110110",
						 "001001100101110100100011",
						 "001001100101110011010000",
						 "001001100101110001111101",
						 "001001100101110000101010",
						 "001001100101101111010111",
						 "001001100101101110000100",
						 "001001100101101100110001",
						 "001001100101101011011110",
						 "001001100101111110111011",
						 "001001100101111101101000",
						 "001001100101111100010101",
						 "001001100101111011000010",
						 "001001100101111001101111",
						 "001001100101111000011100",
						 "001001100101110111001001",
						 "001001100101110101110110",
						 "001001100101110100100011",
						 "001001100101110011010000",
						 "001001100101110001111101",
						 "001001100101110000101010",
						 "001001100101101111010111",
						 "001001100101101110000100",
						 "001001100101101100110001",
						 "001001100101101011011110",
						 "001001100101111110111011",
						 "001001100101111101101000",
						 "001001100101111100010101",
						 "001001100101111011000010",
						 "001001100101111001101111",
						 "001001100101111000011100",
						 "001001100101110111001001",
						 "001001100101110101110110",
						 "001001100101110100100011",
						 "001001100101110011010000",
						 "001001100101110001111101",
						 "001001100101110000101010",
						 "001001100101101111010111",
						 "001001100101101110000100",
						 "001001100101101100110001",
						 "001001100101101011011110",
						 "001001100101111111001010",
						 "001001100101111101110110",
						 "001001100101111100100010",
						 "001001100101111011001110",
						 "001001100101111001111010",
						 "001001100101111000100110",
						 "001001100101110111010010",
						 "001001100101110101111110",
						 "001001100101110100101010",
						 "001001100101110011010110",
						 "001001100101110010000010",
						 "001001100101110000101110",
						 "001001100101101111011010",
						 "001001100101101110000110",
						 "001001100101101100110010",
						 "001001100101101011011110",
						 "001001100101111111001010",
						 "001001100101111101110110",
						 "001001100101111100100010",
						 "001001100101111011001110",
						 "001001100101111001111010",
						 "001001100101111000100110",
						 "001001100101110111010010",
						 "001001100101110101111110",
						 "001001100101110100101010",
						 "001001100101110011010110",
						 "001001100101110010000010",
						 "001001100101110000101110",
						 "001001100101101111011010",
						 "001001100101101110000110",
						 "001001100101101100110010",
						 "001001100101101011011110",
						 "001001100011011100011011",
						 "001001100011011011000110",
						 "001001100011011001110001",
						 "001001100011011000011100",
						 "001001100011010111000111",
						 "001001100011010101110010",
						 "001001100011010100011101",
						 "001001100011010011001000",
						 "001001100011010001110011",
						 "001001100011010000011110",
						 "001001100011001111001001",
						 "001001100011001101110100",
						 "001001100011001100011111",
						 "001001100011001011001010",
						 "001001100011001001110101",
						 "001001100011001000100000",
						 "001001100011011100011011",
						 "001001100011011011000110",
						 "001001100011011001110001",
						 "001001100011011000011100",
						 "001001100011010111000111",
						 "001001100011010101110010",
						 "001001100011010100011101",
						 "001001100011010011001000",
						 "001001100011010001110011",
						 "001001100011010000011110",
						 "001001100011001111001001",
						 "001001100011001101110100",
						 "001001100011001100011111",
						 "001001100011001011001010",
						 "001001100011001001110101",
						 "001001100011001000100000",
						 "001001100011011100011011",
						 "001001100011011011000110",
						 "001001100011011001110001",
						 "001001100011011000011100",
						 "001001100011010111000111",
						 "001001100011010101110010",
						 "001001100011010100011101",
						 "001001100011010011001000",
						 "001001100011010001110011",
						 "001001100011010000011110",
						 "001001100011001111001001",
						 "001001100011001101110100",
						 "001001100011001100011111",
						 "001001100011001011001010",
						 "001001100011001001110101",
						 "001001100011001000100000",
						 "001001100011011100101010",
						 "001001100011011011010100",
						 "001001100011011001111110",
						 "001001100011011000101000",
						 "001001100011010111010010",
						 "001001100011010101111100",
						 "001001100011010100100110",
						 "001001100011010011010000",
						 "001001100011010001111010",
						 "001001100011010000100100",
						 "001001100011001111001110",
						 "001001100011001101111000",
						 "001001100011001100100010",
						 "001001100011001011001100",
						 "001001100011001001110110",
						 "001001100011001000100000",
						 "001001100011011100101010",
						 "001001100011011011010100",
						 "001001100011011001111110",
						 "001001100011011000101000",
						 "001001100011010111010010",
						 "001001100011010101111100",
						 "001001100011010100100110",
						 "001001100011010011010000",
						 "001001100011010001111010",
						 "001001100011010000100100",
						 "001001100011001111001110",
						 "001001100011001101111000",
						 "001001100011001100100010",
						 "001001100011001011001100",
						 "001001100011001001110110",
						 "001001100011001000100000",
						 "001001100011011100101010",
						 "001001100011011011010100",
						 "001001100011011001111110",
						 "001001100011011000101000",
						 "001001100011010111010010",
						 "001001100011010101111100",
						 "001001100011010100100110",
						 "001001100011010011010000",
						 "001001100011010001111010",
						 "001001100011010000100100",
						 "001001100011001111001110",
						 "001001100011001101111000",
						 "001001100011001100100010",
						 "001001100011001011001100",
						 "001001100011001001110110",
						 "001001100011001000100000",
						 "001001100011011100111001",
						 "001001100011011011100010",
						 "001001100011011010001011",
						 "001001100011011000110100",
						 "001001100011010111011101",
						 "001001100011010110000110",
						 "001001100011010100101111",
						 "001001100011010011011000",
						 "001001100011010010000001",
						 "001001100011010000101010",
						 "001001100011001111010011",
						 "001001100011001101111100",
						 "001001100011001100100101",
						 "001001100011001011001110",
						 "001001100011001001110111",
						 "001001100011001000100000",
						 "001001100011011100111001",
						 "001001100011011011100010",
						 "001001100011011010001011",
						 "001001100011011000110100",
						 "001001100011010111011101",
						 "001001100011010110000110",
						 "001001100011010100101111",
						 "001001100011010011011000",
						 "001001100011010010000001",
						 "001001100011010000101010",
						 "001001100011001111010011",
						 "001001100011001101111100",
						 "001001100011001100100101",
						 "001001100011001011001110",
						 "001001100011001001110111",
						 "001001100011001000100000",
						 "001001100000111010001010",
						 "001001100000111000110010",
						 "001001100000110111011010",
						 "001001100000110110000010",
						 "001001100000110100101010",
						 "001001100000110011010010",
						 "001001100000110001111010",
						 "001001100000110000100010",
						 "001001100000101111001010",
						 "001001100000101101110010",
						 "001001100000101100011010",
						 "001001100000101011000010",
						 "001001100000101001101010",
						 "001001100000101000010010",
						 "001001100000100110111010",
						 "001001100000100101100010",
						 "001001100000111010001010",
						 "001001100000111000110010",
						 "001001100000110111011010",
						 "001001100000110110000010",
						 "001001100000110100101010",
						 "001001100000110011010010",
						 "001001100000110001111010",
						 "001001100000110000100010",
						 "001001100000101111001010",
						 "001001100000101101110010",
						 "001001100000101100011010",
						 "001001100000101011000010",
						 "001001100000101001101010",
						 "001001100000101000010010",
						 "001001100000100110111010",
						 "001001100000100101100010",
						 "001001100000111010001010",
						 "001001100000111000110010",
						 "001001100000110111011010",
						 "001001100000110110000010",
						 "001001100000110100101010",
						 "001001100000110011010010",
						 "001001100000110001111010",
						 "001001100000110000100010",
						 "001001100000101111001010",
						 "001001100000101101110010",
						 "001001100000101100011010",
						 "001001100000101011000010",
						 "001001100000101001101010",
						 "001001100000101000010010",
						 "001001100000100110111010",
						 "001001100000100101100010",
						 "001001100000111010011001",
						 "001001100000111001000000",
						 "001001100000110111100111",
						 "001001100000110110001110",
						 "001001100000110100110101",
						 "001001100000110011011100",
						 "001001100000110010000011",
						 "001001100000110000101010",
						 "001001100000101111010001",
						 "001001100000101101111000",
						 "001001100000101100011111",
						 "001001100000101011000110",
						 "001001100000101001101101",
						 "001001100000101000010100",
						 "001001100000100110111011",
						 "001001100000100101100010",
						 "001001100000111010011001",
						 "001001100000111001000000",
						 "001001100000110111100111",
						 "001001100000110110001110",
						 "001001100000110100110101",
						 "001001100000110011011100",
						 "001001100000110010000011",
						 "001001100000110000101010",
						 "001001100000101111010001",
						 "001001100000101101111000",
						 "001001100000101100011111",
						 "001001100000101011000110",
						 "001001100000101001101101",
						 "001001100000101000010100",
						 "001001100000100110111011",
						 "001001100000100101100010",
						 "001001100000111010011001",
						 "001001100000111001000000",
						 "001001100000110111100111",
						 "001001100000110110001110",
						 "001001100000110100110101",
						 "001001100000110011011100",
						 "001001100000110010000011",
						 "001001100000110000101010",
						 "001001100000101111010001",
						 "001001100000101101111000",
						 "001001100000101100011111",
						 "001001100000101011000110",
						 "001001100000101001101101",
						 "001001100000101000010100",
						 "001001100000100110111011",
						 "001001100000100101100010",
						 "001001100000111010101000",
						 "001001100000111001001110",
						 "001001100000110111110100",
						 "001001100000110110011010",
						 "001001100000110101000000",
						 "001001100000110011100110",
						 "001001100000110010001100",
						 "001001100000110000110010",
						 "001001100000101111011000",
						 "001001100000101101111110",
						 "001001100000101100100100",
						 "001001100000101011001010",
						 "001001100000101001110000",
						 "001001100000101000010110",
						 "001001100000100110111100",
						 "001001100000100101100010",
						 "001001011110010111101010",
						 "001001011110010110010000",
						 "001001011110010100110110",
						 "001001011110010011011100",
						 "001001011110010010000010",
						 "001001011110010000101000",
						 "001001011110001111001110",
						 "001001011110001101110100",
						 "001001011110001100011010",
						 "001001011110001011000000",
						 "001001011110001001100110",
						 "001001011110001000001100",
						 "001001011110000110110010",
						 "001001011110000101011000",
						 "001001011110000011111110",
						 "001001011110000010100100",
						 "001001011110010111101010",
						 "001001011110010110010000",
						 "001001011110010100110110",
						 "001001011110010011011100",
						 "001001011110010010000010",
						 "001001011110010000101000",
						 "001001011110001111001110",
						 "001001011110001101110100",
						 "001001011110001100011010",
						 "001001011110001011000000",
						 "001001011110001001100110",
						 "001001011110001000001100",
						 "001001011110000110110010",
						 "001001011110000101011000",
						 "001001011110000011111110",
						 "001001011110000010100100",
						 "001001011110010111111001",
						 "001001011110010110011110",
						 "001001011110010101000011",
						 "001001011110010011101000",
						 "001001011110010010001101",
						 "001001011110010000110010",
						 "001001011110001111010111",
						 "001001011110001101111100",
						 "001001011110001100100001",
						 "001001011110001011000110",
						 "001001011110001001101011",
						 "001001011110001000010000",
						 "001001011110000110110101",
						 "001001011110000101011010",
						 "001001011110000011111111",
						 "001001011110000010100100",
						 "001001011110010111111001",
						 "001001011110010110011110",
						 "001001011110010101000011",
						 "001001011110010011101000",
						 "001001011110010010001101",
						 "001001011110010000110010",
						 "001001011110001111010111",
						 "001001011110001101111100",
						 "001001011110001100100001",
						 "001001011110001011000110",
						 "001001011110001001101011",
						 "001001011110001000010000",
						 "001001011110000110110101",
						 "001001011110000101011010",
						 "001001011110000011111111",
						 "001001011110000010100100",
						 "001001011110011000001000",
						 "001001011110010110101100",
						 "001001011110010101010000",
						 "001001011110010011110100",
						 "001001011110010010011000",
						 "001001011110010000111100",
						 "001001011110001111100000",
						 "001001011110001110000100",
						 "001001011110001100101000",
						 "001001011110001011001100",
						 "001001011110001001110000",
						 "001001011110001000010100",
						 "001001011110000110111000",
						 "001001011110000101011100",
						 "001001011110000100000000",
						 "001001011110000010100100",
						 "001001011110011000001000",
						 "001001011110010110101100",
						 "001001011110010101010000",
						 "001001011110010011110100",
						 "001001011110010010011000",
						 "001001011110010000111100",
						 "001001011110001111100000",
						 "001001011110001110000100",
						 "001001011110001100101000",
						 "001001011110001011001100",
						 "001001011110001001110000",
						 "001001011110001000010100",
						 "001001011110000110111000",
						 "001001011110000101011100",
						 "001001011110000100000000",
						 "001001011110000010100100",
						 "001001011110011000001000",
						 "001001011110010110101100",
						 "001001011110010101010000",
						 "001001011110010011110100",
						 "001001011110010010011000",
						 "001001011110010000111100",
						 "001001011110001111100000",
						 "001001011110001110000100",
						 "001001011110001100101000",
						 "001001011110001011001100",
						 "001001011110001001110000",
						 "001001011110001000010100",
						 "001001011110000110111000",
						 "001001011110000101011100",
						 "001001011110000100000000",
						 "001001011110000010100100",
						 "001001011011110101011001",
						 "001001011011110011111100",
						 "001001011011110010011111",
						 "001001011011110001000010",
						 "001001011011101111100101",
						 "001001011011101110001000",
						 "001001011011101100101011",
						 "001001011011101011001110",
						 "001001011011101001110001",
						 "001001011011101000010100",
						 "001001011011100110110111",
						 "001001011011100101011010",
						 "001001011011100011111101",
						 "001001011011100010100000",
						 "001001011011100001000011",
						 "001001011011011111100110",
						 "001001011011110101011001",
						 "001001011011110011111100",
						 "001001011011110010011111",
						 "001001011011110001000010",
						 "001001011011101111100101",
						 "001001011011101110001000",
						 "001001011011101100101011",
						 "001001011011101011001110",
						 "001001011011101001110001",
						 "001001011011101000010100",
						 "001001011011100110110111",
						 "001001011011100101011010",
						 "001001011011100011111101",
						 "001001011011100010100000",
						 "001001011011100001000011",
						 "001001011011011111100110",
						 "001001011011110101011001",
						 "001001011011110011111100",
						 "001001011011110010011111",
						 "001001011011110001000010",
						 "001001011011101111100101",
						 "001001011011101110001000",
						 "001001011011101100101011",
						 "001001011011101011001110",
						 "001001011011101001110001",
						 "001001011011101000010100",
						 "001001011011100110110111",
						 "001001011011100101011010",
						 "001001011011100011111101",
						 "001001011011100010100000",
						 "001001011011100001000011",
						 "001001011011011111100110",
						 "001001011011110101101000",
						 "001001011011110100001010",
						 "001001011011110010101100",
						 "001001011011110001001110",
						 "001001011011101111110000",
						 "001001011011101110010010",
						 "001001011011101100110100",
						 "001001011011101011010110",
						 "001001011011101001111000",
						 "001001011011101000011010",
						 "001001011011100110111100",
						 "001001011011100101011110",
						 "001001011011100100000000",
						 "001001011011100010100010",
						 "001001011011100001000100",
						 "001001011011011111100110",
						 "001001011011110101101000",
						 "001001011011110100001010",
						 "001001011011110010101100",
						 "001001011011110001001110",
						 "001001011011101111110000",
						 "001001011011101110010010",
						 "001001011011101100110100",
						 "001001011011101011010110",
						 "001001011011101001111000",
						 "001001011011101000011010",
						 "001001011011100110111100",
						 "001001011011100101011110",
						 "001001011011100100000000",
						 "001001011011100010100010",
						 "001001011011100001000100",
						 "001001011011011111100110",
						 "001001011011110101101000",
						 "001001011011110100001010",
						 "001001011011110010101100",
						 "001001011011110001001110",
						 "001001011011101111110000",
						 "001001011011101110010010",
						 "001001011011101100110100",
						 "001001011011101011010110",
						 "001001011011101001111000",
						 "001001011011101000011010",
						 "001001011011100110111100",
						 "001001011011100101011110",
						 "001001011011100100000000",
						 "001001011011100010100010",
						 "001001011011100001000100",
						 "001001011011011111100110",
						 "001001011011110101110111",
						 "001001011011110100011000",
						 "001001011011110010111001",
						 "001001011011110001011010",
						 "001001011011101111111011",
						 "001001011011101110011100",
						 "001001011011101100111101",
						 "001001011011101011011110",
						 "001001011011101001111111",
						 "001001011011101000100000",
						 "001001011011100111000001",
						 "001001011011100101100010",
						 "001001011011100100000011",
						 "001001011011100010100100",
						 "001001011011100001000101",
						 "001001011011011111100110",
						 "001001011001010010111001",
						 "001001011001010001011010",
						 "001001011001001111111011",
						 "001001011001001110011100",
						 "001001011001001100111101",
						 "001001011001001011011110",
						 "001001011001001001111111",
						 "001001011001001000100000",
						 "001001011001000111000001",
						 "001001011001000101100010",
						 "001001011001000100000011",
						 "001001011001000010100100",
						 "001001011001000001000101",
						 "001001011000111111100110",
						 "001001011000111110000111",
						 "001001011000111100101000",
						 "001001011001010011001000",
						 "001001011001010001101000",
						 "001001011001010000001000",
						 "001001011001001110101000",
						 "001001011001001101001000",
						 "001001011001001011101000",
						 "001001011001001010001000",
						 "001001011001001000101000",
						 "001001011001000111001000",
						 "001001011001000101101000",
						 "001001011001000100001000",
						 "001001011001000010101000",
						 "001001011001000001001000",
						 "001001011000111111101000",
						 "001001011000111110001000",
						 "001001011000111100101000",
						 "001001011001010011001000",
						 "001001011001010001101000",
						 "001001011001010000001000",
						 "001001011001001110101000",
						 "001001011001001101001000",
						 "001001011001001011101000",
						 "001001011001001010001000",
						 "001001011001001000101000",
						 "001001011001000111001000",
						 "001001011001000101101000",
						 "001001011001000100001000",
						 "001001011001000010101000",
						 "001001011001000001001000",
						 "001001011000111111101000",
						 "001001011000111110001000",
						 "001001011000111100101000",
						 "001001011001010011001000",
						 "001001011001010001101000",
						 "001001011001010000001000",
						 "001001011001001110101000",
						 "001001011001001101001000",
						 "001001011001001011101000",
						 "001001011001001010001000",
						 "001001011001001000101000",
						 "001001011001000111001000",
						 "001001011001000101101000",
						 "001001011001000100001000",
						 "001001011001000010101000",
						 "001001011001000001001000",
						 "001001011000111111101000",
						 "001001011000111110001000",
						 "001001011000111100101000",
						 "001001011001010011010111",
						 "001001011001010001110110",
						 "001001011001010000010101",
						 "001001011001001110110100",
						 "001001011001001101010011",
						 "001001011001001011110010",
						 "001001011001001010010001",
						 "001001011001001000110000",
						 "001001011001000111001111",
						 "001001011001000101101110",
						 "001001011001000100001101",
						 "001001011001000010101100",
						 "001001011001000001001011",
						 "001001011000111111101010",
						 "001001011000111110001001",
						 "001001011000111100101000",
						 "001001011001010011010111",
						 "001001011001010001110110",
						 "001001011001010000010101",
						 "001001011001001110110100",
						 "001001011001001101010011",
						 "001001011001001011110010",
						 "001001011001001010010001",
						 "001001011001001000110000",
						 "001001011001000111001111",
						 "001001011001000101101110",
						 "001001011001000100001101",
						 "001001011001000010101100",
						 "001001011001000001001011",
						 "001001011000111111101010",
						 "001001011000111110001001",
						 "001001011000111100101000",
						 "001001011001010011010111",
						 "001001011001010001110110",
						 "001001011001010000010101",
						 "001001011001001110110100",
						 "001001011001001101010011",
						 "001001011001001011110010",
						 "001001011001001010010001",
						 "001001011001001000110000",
						 "001001011001000111001111",
						 "001001011001000101101110",
						 "001001011001000100001101",
						 "001001011001000010101100",
						 "001001011001000001001011",
						 "001001011000111111101010",
						 "001001011000111110001001",
						 "001001011000111100101000",
						 "001001010110110000101000",
						 "001001010110101111000110",
						 "001001010110101101100100",
						 "001001010110101100000010",
						 "001001010110101010100000",
						 "001001010110101000111110",
						 "001001010110100111011100",
						 "001001010110100101111010",
						 "001001010110100100011000",
						 "001001010110100010110110",
						 "001001010110100001010100",
						 "001001010110011111110010",
						 "001001010110011110010000",
						 "001001010110011100101110",
						 "001001010110011011001100",
						 "001001010110011001101010",
						 "001001010110110000101000",
						 "001001010110101111000110",
						 "001001010110101101100100",
						 "001001010110101100000010",
						 "001001010110101010100000",
						 "001001010110101000111110",
						 "001001010110100111011100",
						 "001001010110100101111010",
						 "001001010110100100011000",
						 "001001010110100010110110",
						 "001001010110100001010100",
						 "001001010110011111110010",
						 "001001010110011110010000",
						 "001001010110011100101110",
						 "001001010110011011001100",
						 "001001010110011001101010",
						 "001001010110110000101000",
						 "001001010110101111000110",
						 "001001010110101101100100",
						 "001001010110101100000010",
						 "001001010110101010100000",
						 "001001010110101000111110",
						 "001001010110100111011100",
						 "001001010110100101111010",
						 "001001010110100100011000",
						 "001001010110100010110110",
						 "001001010110100001010100",
						 "001001010110011111110010",
						 "001001010110011110010000",
						 "001001010110011100101110",
						 "001001010110011011001100",
						 "001001010110011001101010",
						 "001001010110110000110111",
						 "001001010110101111010100",
						 "001001010110101101110001",
						 "001001010110101100001110",
						 "001001010110101010101011",
						 "001001010110101001001000",
						 "001001010110100111100101",
						 "001001010110100110000010",
						 "001001010110100100011111",
						 "001001010110100010111100",
						 "001001010110100001011001",
						 "001001010110011111110110",
						 "001001010110011110010011",
						 "001001010110011100110000",
						 "001001010110011011001101",
						 "001001010110011001101010",
						 "001001010110110000110111",
						 "001001010110101111010100",
						 "001001010110101101110001",
						 "001001010110101100001110",
						 "001001010110101010101011",
						 "001001010110101001001000",
						 "001001010110100111100101",
						 "001001010110100110000010",
						 "001001010110100100011111",
						 "001001010110100010111100",
						 "001001010110100001011001",
						 "001001010110011111110110",
						 "001001010110011110010011",
						 "001001010110011100110000",
						 "001001010110011011001101",
						 "001001010110011001101010",
						 "001001010110110001000110",
						 "001001010110101111100010",
						 "001001010110101101111110",
						 "001001010110101100011010",
						 "001001010110101010110110",
						 "001001010110101001010010",
						 "001001010110100111101110",
						 "001001010110100110001010",
						 "001001010110100100100110",
						 "001001010110100011000010",
						 "001001010110100001011110",
						 "001001010110011111111010",
						 "001001010110011110010110",
						 "001001010110011100110010",
						 "001001010110011011001110",
						 "001001010110011001101010",
						 "001001010110110001000110",
						 "001001010110101111100010",
						 "001001010110101101111110",
						 "001001010110101100011010",
						 "001001010110101010110110",
						 "001001010110101001010010",
						 "001001010110100111101110",
						 "001001010110100110001010",
						 "001001010110100100100110",
						 "001001010110100011000010",
						 "001001010110100001011110",
						 "001001010110011111111010",
						 "001001010110011110010110",
						 "001001010110011100110010",
						 "001001010110011011001110",
						 "001001010110011001101010",
						 "001001010100001110001000",
						 "001001010100001100100100",
						 "001001010100001011000000",
						 "001001010100001001011100",
						 "001001010100000111111000",
						 "001001010100000110010100",
						 "001001010100000100110000",
						 "001001010100000011001100",
						 "001001010100000001101000",
						 "001001010100000000000100",
						 "001001010011111110100000",
						 "001001010011111100111100",
						 "001001010011111011011000",
						 "001001010011111001110100",
						 "001001010011111000010000",
						 "001001010011110110101100",
						 "001001010100001110010111",
						 "001001010100001100110010",
						 "001001010100001011001101",
						 "001001010100001001101000",
						 "001001010100001000000011",
						 "001001010100000110011110",
						 "001001010100000100111001",
						 "001001010100000011010100",
						 "001001010100000001101111",
						 "001001010100000000001010",
						 "001001010011111110100101",
						 "001001010011111101000000",
						 "001001010011111011011011",
						 "001001010011111001110110",
						 "001001010011111000010001",
						 "001001010011110110101100",
						 "001001010100001110010111",
						 "001001010100001100110010",
						 "001001010100001011001101",
						 "001001010100001001101000",
						 "001001010100001000000011",
						 "001001010100000110011110",
						 "001001010100000100111001",
						 "001001010100000011010100",
						 "001001010100000001101111",
						 "001001010100000000001010",
						 "001001010011111110100101",
						 "001001010011111101000000",
						 "001001010011111011011011",
						 "001001010011111001110110",
						 "001001010011111000010001",
						 "001001010011110110101100",
						 "001001010100001110010111",
						 "001001010100001100110010",
						 "001001010100001011001101",
						 "001001010100001001101000",
						 "001001010100001000000011",
						 "001001010100000110011110",
						 "001001010100000100111001",
						 "001001010100000011010100",
						 "001001010100000001101111",
						 "001001010100000000001010",
						 "001001010011111110100101",
						 "001001010011111101000000",
						 "001001010011111011011011",
						 "001001010011111001110110",
						 "001001010011111000010001",
						 "001001010011110110101100",
						 "001001010100001110100110",
						 "001001010100001101000000",
						 "001001010100001011011010",
						 "001001010100001001110100",
						 "001001010100001000001110",
						 "001001010100000110101000",
						 "001001010100000101000010",
						 "001001010100000011011100",
						 "001001010100000001110110",
						 "001001010100000000010000",
						 "001001010011111110101010",
						 "001001010011111101000100",
						 "001001010011111011011110",
						 "001001010011111001111000",
						 "001001010011111000010010",
						 "001001010011110110101100",
						 "001001010100001110100110",
						 "001001010100001101000000",
						 "001001010100001011011010",
						 "001001010100001001110100",
						 "001001010100001000001110",
						 "001001010100000110101000",
						 "001001010100000101000010",
						 "001001010100000011011100",
						 "001001010100000001110110",
						 "001001010100000000010000",
						 "001001010011111110101010",
						 "001001010011111101000100",
						 "001001010011111011011110",
						 "001001010011111001111000",
						 "001001010011111000010010",
						 "001001010011110110101100",
						 "001001010001101011101000",
						 "001001010001101010000010",
						 "001001010001101000011100",
						 "001001010001100110110110",
						 "001001010001100101010000",
						 "001001010001100011101010",
						 "001001010001100010000100",
						 "001001010001100000011110",
						 "001001010001011110111000",
						 "001001010001011101010010",
						 "001001010001011011101100",
						 "001001010001011010000110",
						 "001001010001011000100000",
						 "001001010001010110111010",
						 "001001010001010101010100",
						 "001001010001010011101110",
						 "001001010001101011110111",
						 "001001010001101010010000",
						 "001001010001101000101001",
						 "001001010001100111000010",
						 "001001010001100101011011",
						 "001001010001100011110100",
						 "001001010001100010001101",
						 "001001010001100000100110",
						 "001001010001011110111111",
						 "001001010001011101011000",
						 "001001010001011011110001",
						 "001001010001011010001010",
						 "001001010001011000100011",
						 "001001010001010110111100",
						 "001001010001010101010101",
						 "001001010001010011101110",
						 "001001010001101011110111",
						 "001001010001101010010000",
						 "001001010001101000101001",
						 "001001010001100111000010",
						 "001001010001100101011011",
						 "001001010001100011110100",
						 "001001010001100010001101",
						 "001001010001100000100110",
						 "001001010001011110111111",
						 "001001010001011101011000",
						 "001001010001011011110001",
						 "001001010001011010001010",
						 "001001010001011000100011",
						 "001001010001010110111100",
						 "001001010001010101010101",
						 "001001010001010011101110",
						 "001001010001101100000110",
						 "001001010001101010011110",
						 "001001010001101000110110",
						 "001001010001100111001110",
						 "001001010001100101100110",
						 "001001010001100011111110",
						 "001001010001100010010110",
						 "001001010001100000101110",
						 "001001010001011111000110",
						 "001001010001011101011110",
						 "001001010001011011110110",
						 "001001010001011010001110",
						 "001001010001011000100110",
						 "001001010001010110111110",
						 "001001010001010101010110",
						 "001001010001010011101110",
						 "001001010001101100000110",
						 "001001010001101010011110",
						 "001001010001101000110110",
						 "001001010001100111001110",
						 "001001010001100101100110",
						 "001001010001100011111110",
						 "001001010001100010010110",
						 "001001010001100000101110",
						 "001001010001011111000110",
						 "001001010001011101011110",
						 "001001010001011011110110",
						 "001001010001011010001110",
						 "001001010001011000100110",
						 "001001010001010110111110",
						 "001001010001010101010110",
						 "001001010001010011101110",
						 "001001010001101100000110",
						 "001001010001101010011110",
						 "001001010001101000110110",
						 "001001010001100111001110",
						 "001001010001100101100110",
						 "001001010001100011111110",
						 "001001010001100010010110",
						 "001001010001100000101110",
						 "001001010001011111000110",
						 "001001010001011101011110",
						 "001001010001011011110110",
						 "001001010001011010001110",
						 "001001010001011000100110",
						 "001001010001010110111110",
						 "001001010001010101010110",
						 "001001010001010011101110",
						 "001001001111001001010111",
						 "001001001111000111101110",
						 "001001001111000110000101",
						 "001001001111000100011100",
						 "001001001111000010110011",
						 "001001001111000001001010",
						 "001001001110111111100001",
						 "001001001110111101111000",
						 "001001001110111100001111",
						 "001001001110111010100110",
						 "001001001110111000111101",
						 "001001001110110111010100",
						 "001001001110110101101011",
						 "001001001110110100000010",
						 "001001001110110010011001",
						 "001001001110110000110000",
						 "001001001111001001010111",
						 "001001001111000111101110",
						 "001001001111000110000101",
						 "001001001111000100011100",
						 "001001001111000010110011",
						 "001001001111000001001010",
						 "001001001110111111100001",
						 "001001001110111101111000",
						 "001001001110111100001111",
						 "001001001110111010100110",
						 "001001001110111000111101",
						 "001001001110110111010100",
						 "001001001110110101101011",
						 "001001001110110100000010",
						 "001001001110110010011001",
						 "001001001110110000110000",
						 "001001001111001001010111",
						 "001001001111000111101110",
						 "001001001111000110000101",
						 "001001001111000100011100",
						 "001001001111000010110011",
						 "001001001111000001001010",
						 "001001001110111111100001",
						 "001001001110111101111000",
						 "001001001110111100001111",
						 "001001001110111010100110",
						 "001001001110111000111101",
						 "001001001110110111010100",
						 "001001001110110101101011",
						 "001001001110110100000010",
						 "001001001110110010011001",
						 "001001001110110000110000",
						 "001001001111001001100110",
						 "001001001111000111111100",
						 "001001001111000110010010",
						 "001001001111000100101000",
						 "001001001111000010111110",
						 "001001001111000001010100",
						 "001001001110111111101010",
						 "001001001110111110000000",
						 "001001001110111100010110",
						 "001001001110111010101100",
						 "001001001110111001000010",
						 "001001001110110111011000",
						 "001001001110110101101110",
						 "001001001110110100000100",
						 "001001001110110010011010",
						 "001001001110110000110000",
						 "001001001111001001100110",
						 "001001001111000111111100",
						 "001001001111000110010010",
						 "001001001111000100101000",
						 "001001001111000010111110",
						 "001001001111000001010100",
						 "001001001110111111101010",
						 "001001001110111110000000",
						 "001001001110111100010110",
						 "001001001110111010101100",
						 "001001001110111001000010",
						 "001001001110110111011000",
						 "001001001110110101101110",
						 "001001001110110100000100",
						 "001001001110110010011010",
						 "001001001110110000110000",
						 "001001001111001001100110",
						 "001001001111000111111100",
						 "001001001111000110010010",
						 "001001001111000100101000",
						 "001001001111000010111110",
						 "001001001111000001010100",
						 "001001001110111111101010",
						 "001001001110111110000000",
						 "001001001110111100010110",
						 "001001001110111010101100",
						 "001001001110111001000010",
						 "001001001110110111011000",
						 "001001001110110101101110",
						 "001001001110110100000100",
						 "001001001110110010011010",
						 "001001001110110000110000",
						 "001001001111001001110101",
						 "001001001111001000001010",
						 "001001001111000110011111",
						 "001001001111000100110100",
						 "001001001111000011001001",
						 "001001001111000001011110",
						 "001001001110111111110011",
						 "001001001110111110001000",
						 "001001001110111100011101",
						 "001001001110111010110010",
						 "001001001110111001000111",
						 "001001001110110111011100",
						 "001001001110110101110001",
						 "001001001110110100000110",
						 "001001001110110010011011",
						 "001001001110110000110000",
						 "001001001100100110110111",
						 "001001001100100101001100",
						 "001001001100100011100001",
						 "001001001100100001110110",
						 "001001001100100000001011",
						 "001001001100011110100000",
						 "001001001100011100110101",
						 "001001001100011011001010",
						 "001001001100011001011111",
						 "001001001100010111110100",
						 "001001001100010110001001",
						 "001001001100010100011110",
						 "001001001100010010110011",
						 "001001001100010001001000",
						 "001001001100001111011101",
						 "001001001100001101110010",
						 "001001001100100110110111",
						 "001001001100100101001100",
						 "001001001100100011100001",
						 "001001001100100001110110",
						 "001001001100100000001011",
						 "001001001100011110100000",
						 "001001001100011100110101",
						 "001001001100011011001010",
						 "001001001100011001011111",
						 "001001001100010111110100",
						 "001001001100010110001001",
						 "001001001100010100011110",
						 "001001001100010010110011",
						 "001001001100010001001000",
						 "001001001100001111011101",
						 "001001001100001101110010",
						 "001001001100100111000110",
						 "001001001100100101011010",
						 "001001001100100011101110",
						 "001001001100100010000010",
						 "001001001100100000010110",
						 "001001001100011110101010",
						 "001001001100011100111110",
						 "001001001100011011010010",
						 "001001001100011001100110",
						 "001001001100010111111010",
						 "001001001100010110001110",
						 "001001001100010100100010",
						 "001001001100010010110110",
						 "001001001100010001001010",
						 "001001001100001111011110",
						 "001001001100001101110010",
						 "001001001100100111000110",
						 "001001001100100101011010",
						 "001001001100100011101110",
						 "001001001100100010000010",
						 "001001001100100000010110",
						 "001001001100011110101010",
						 "001001001100011100111110",
						 "001001001100011011010010",
						 "001001001100011001100110",
						 "001001001100010111111010",
						 "001001001100010110001110",
						 "001001001100010100100010",
						 "001001001100010010110110",
						 "001001001100010001001010",
						 "001001001100001111011110",
						 "001001001100001101110010",
						 "001001001100100111000110",
						 "001001001100100101011010",
						 "001001001100100011101110",
						 "001001001100100010000010",
						 "001001001100100000010110",
						 "001001001100011110101010",
						 "001001001100011100111110",
						 "001001001100011011010010",
						 "001001001100011001100110",
						 "001001001100010111111010",
						 "001001001100010110001110",
						 "001001001100010100100010",
						 "001001001100010010110110",
						 "001001001100010001001010",
						 "001001001100001111011110",
						 "001001001100001101110010",
						 "001001001100100111010101",
						 "001001001100100101101000",
						 "001001001100100011111011",
						 "001001001100100010001110",
						 "001001001100100000100001",
						 "001001001100011110110100",
						 "001001001100011101000111",
						 "001001001100011011011010",
						 "001001001100011001101101",
						 "001001001100011000000000",
						 "001001001100010110010011",
						 "001001001100010100100110",
						 "001001001100010010111001",
						 "001001001100010001001100",
						 "001001001100001111011111",
						 "001001001100001101110010",
						 "001001001010000100010111",
						 "001001001010000010101010",
						 "001001001010000000111101",
						 "001001001001111111010000",
						 "001001001001111101100011",
						 "001001001001111011110110",
						 "001001001001111010001001",
						 "001001001001111000011100",
						 "001001001001110110101111",
						 "001001001001110101000010",
						 "001001001001110011010101",
						 "001001001001110001101000",
						 "001001001001101111111011",
						 "001001001001101110001110",
						 "001001001001101100100001",
						 "001001001001101010110100",
						 "001001001010000100100110",
						 "001001001010000010111000",
						 "001001001010000001001010",
						 "001001001001111111011100",
						 "001001001001111101101110",
						 "001001001001111100000000",
						 "001001001001111010010010",
						 "001001001001111000100100",
						 "001001001001110110110110",
						 "001001001001110101001000",
						 "001001001001110011011010",
						 "001001001001110001101100",
						 "001001001001101111111110",
						 "001001001001101110010000",
						 "001001001001101100100010",
						 "001001001001101010110100",
						 "001001001010000100100110",
						 "001001001010000010111000",
						 "001001001010000001001010",
						 "001001001001111111011100",
						 "001001001001111101101110",
						 "001001001001111100000000",
						 "001001001001111010010010",
						 "001001001001111000100100",
						 "001001001001110110110110",
						 "001001001001110101001000",
						 "001001001001110011011010",
						 "001001001001110001101100",
						 "001001001001101111111110",
						 "001001001001101110010000",
						 "001001001001101100100010",
						 "001001001001101010110100",
						 "001001001010000100100110",
						 "001001001010000010111000",
						 "001001001010000001001010",
						 "001001001001111111011100",
						 "001001001001111101101110",
						 "001001001001111100000000",
						 "001001001001111010010010",
						 "001001001001111000100100",
						 "001001001001110110110110",
						 "001001001001110101001000",
						 "001001001001110011011010",
						 "001001001001110001101100",
						 "001001001001101111111110",
						 "001001001001101110010000",
						 "001001001001101100100010",
						 "001001001001101010110100",
						 "001001001010000100110101",
						 "001001001010000011000110",
						 "001001001010000001010111",
						 "001001001001111111101000",
						 "001001001001111101111001",
						 "001001001001111100001010",
						 "001001001001111010011011",
						 "001001001001111000101100",
						 "001001001001110110111101",
						 "001001001001110101001110",
						 "001001001001110011011111",
						 "001001001001110001110000",
						 "001001001001110000000001",
						 "001001001001101110010010",
						 "001001001001101100100011",
						 "001001001001101010110100",
						 "001001001010000100110101",
						 "001001001010000011000110",
						 "001001001010000001010111",
						 "001001001001111111101000",
						 "001001001001111101111001",
						 "001001001001111100001010",
						 "001001001001111010011011",
						 "001001001001111000101100",
						 "001001001001110110111101",
						 "001001001001110101001110",
						 "001001001001110011011111",
						 "001001001001110001110000",
						 "001001001001110000000001",
						 "001001001001101110010010",
						 "001001001001101100100011",
						 "001001001001101010110100",
						 "001001000111100001110111",
						 "001001000111100000001000",
						 "001001000111011110011001",
						 "001001000111011100101010",
						 "001001000111011010111011",
						 "001001000111011001001100",
						 "001001000111010111011101",
						 "001001000111010101101110",
						 "001001000111010011111111",
						 "001001000111010010010000",
						 "001001000111010000100001",
						 "001001000111001110110010",
						 "001001000111001101000011",
						 "001001000111001011010100",
						 "001001000111001001100101",
						 "001001000111000111110110",
						 "001001000111100010000110",
						 "001001000111100000010110",
						 "001001000111011110100110",
						 "001001000111011100110110",
						 "001001000111011011000110",
						 "001001000111011001010110",
						 "001001000111010111100110",
						 "001001000111010101110110",
						 "001001000111010100000110",
						 "001001000111010010010110",
						 "001001000111010000100110",
						 "001001000111001110110110",
						 "001001000111001101000110",
						 "001001000111001011010110",
						 "001001000111001001100110",
						 "001001000111000111110110",
						 "001001000111100010000110",
						 "001001000111100000010110",
						 "001001000111011110100110",
						 "001001000111011100110110",
						 "001001000111011011000110",
						 "001001000111011001010110",
						 "001001000111010111100110",
						 "001001000111010101110110",
						 "001001000111010100000110",
						 "001001000111010010010110",
						 "001001000111010000100110",
						 "001001000111001110110110",
						 "001001000111001101000110",
						 "001001000111001011010110",
						 "001001000111001001100110",
						 "001001000111000111110110",
						 "001001000111100010000110",
						 "001001000111100000010110",
						 "001001000111011110100110",
						 "001001000111011100110110",
						 "001001000111011011000110",
						 "001001000111011001010110",
						 "001001000111010111100110",
						 "001001000111010101110110",
						 "001001000111010100000110",
						 "001001000111010010010110",
						 "001001000111010000100110",
						 "001001000111001110110110",
						 "001001000111001101000110",
						 "001001000111001011010110",
						 "001001000111001001100110",
						 "001001000111000111110110",
						 "001001000111100010010101",
						 "001001000111100000100100",
						 "001001000111011110110011",
						 "001001000111011101000010",
						 "001001000111011011010001",
						 "001001000111011001100000",
						 "001001000111010111101111",
						 "001001000111010101111110",
						 "001001000111010100001101",
						 "001001000111010010011100",
						 "001001000111010000101011",
						 "001001000111001110111010",
						 "001001000111001101001001",
						 "001001000111001011011000",
						 "001001000111001001100111",
						 "001001000111000111110110",
						 "001001000100111111010111",
						 "001001000100111101100110",
						 "001001000100111011110101",
						 "001001000100111010000100",
						 "001001000100111000010011",
						 "001001000100110110100010",
						 "001001000100110100110001",
						 "001001000100110011000000",
						 "001001000100110001001111",
						 "001001000100101111011110",
						 "001001000100101101101101",
						 "001001000100101011111100",
						 "001001000100101010001011",
						 "001001000100101000011010",
						 "001001000100100110101001",
						 "001001000100100100111000",
						 "001001000100111111010111",
						 "001001000100111101100110",
						 "001001000100111011110101",
						 "001001000100111010000100",
						 "001001000100111000010011",
						 "001001000100110110100010",
						 "001001000100110100110001",
						 "001001000100110011000000",
						 "001001000100110001001111",
						 "001001000100101111011110",
						 "001001000100101101101101",
						 "001001000100101011111100",
						 "001001000100101010001011",
						 "001001000100101000011010",
						 "001001000100100110101001",
						 "001001000100100100111000",
						 "001001000100111111100110",
						 "001001000100111101110100",
						 "001001000100111100000010",
						 "001001000100111010010000",
						 "001001000100111000011110",
						 "001001000100110110101100",
						 "001001000100110100111010",
						 "001001000100110011001000",
						 "001001000100110001010110",
						 "001001000100101111100100",
						 "001001000100101101110010",
						 "001001000100101100000000",
						 "001001000100101010001110",
						 "001001000100101000011100",
						 "001001000100100110101010",
						 "001001000100100100111000",
						 "001001000100111111100110",
						 "001001000100111101110100",
						 "001001000100111100000010",
						 "001001000100111010010000",
						 "001001000100111000011110",
						 "001001000100110110101100",
						 "001001000100110100111010",
						 "001001000100110011001000",
						 "001001000100110001010110",
						 "001001000100101111100100",
						 "001001000100101101110010",
						 "001001000100101100000000",
						 "001001000100101010001110",
						 "001001000100101000011100",
						 "001001000100100110101010",
						 "001001000100100100111000",
						 "001001000100111111100110",
						 "001001000100111101110100",
						 "001001000100111100000010",
						 "001001000100111010010000",
						 "001001000100111000011110",
						 "001001000100110110101100",
						 "001001000100110100111010",
						 "001001000100110011001000",
						 "001001000100110001010110",
						 "001001000100101111100100",
						 "001001000100101101110010",
						 "001001000100101100000000",
						 "001001000100101010001110",
						 "001001000100101000011100",
						 "001001000100100110101010",
						 "001001000100100100111000",
						 "001001000100111111110101",
						 "001001000100111110000010",
						 "001001000100111100001111",
						 "001001000100111010011100",
						 "001001000100111000101001",
						 "001001000100110110110110",
						 "001001000100110101000011",
						 "001001000100110011010000",
						 "001001000100110001011101",
						 "001001000100101111101010",
						 "001001000100101101110111",
						 "001001000100101100000100",
						 "001001000100101010010001",
						 "001001000100101000011110",
						 "001001000100100110101011",
						 "001001000100100100111000",
						 "001001000010011100110111",
						 "001001000010011011000100",
						 "001001000010011001010001",
						 "001001000010010111011110",
						 "001001000010010101101011",
						 "001001000010010011111000",
						 "001001000010010010000101",
						 "001001000010010000010010",
						 "001001000010001110011111",
						 "001001000010001100101100",
						 "001001000010001010111001",
						 "001001000010001001000110",
						 "001001000010000111010011",
						 "001001000010000101100000",
						 "001001000010000011101101",
						 "001001000010000001111010",
						 "001001000010011101000110",
						 "001001000010011011010010",
						 "001001000010011001011110",
						 "001001000010010111101010",
						 "001001000010010101110110",
						 "001001000010010100000010",
						 "001001000010010010001110",
						 "001001000010010000011010",
						 "001001000010001110100110",
						 "001001000010001100110010",
						 "001001000010001010111110",
						 "001001000010001001001010",
						 "001001000010000111010110",
						 "001001000010000101100010",
						 "001001000010000011101110",
						 "001001000010000001111010",
						 "001001000010011101000110",
						 "001001000010011011010010",
						 "001001000010011001011110",
						 "001001000010010111101010",
						 "001001000010010101110110",
						 "001001000010010100000010",
						 "001001000010010010001110",
						 "001001000010010000011010",
						 "001001000010001110100110",
						 "001001000010001100110010",
						 "001001000010001010111110",
						 "001001000010001001001010",
						 "001001000010000111010110",
						 "001001000010000101100010",
						 "001001000010000011101110",
						 "001001000010000001111010",
						 "001001000010011101000110",
						 "001001000010011011010010",
						 "001001000010011001011110",
						 "001001000010010111101010",
						 "001001000010010101110110",
						 "001001000010010100000010",
						 "001001000010010010001110",
						 "001001000010010000011010",
						 "001001000010001110100110",
						 "001001000010001100110010",
						 "001001000010001010111110",
						 "001001000010001001001010",
						 "001001000010000111010110",
						 "001001000010000101100010",
						 "001001000010000011101110",
						 "001001000010000001111010",
						 "001001000010011101010101",
						 "001001000010011011100000",
						 "001001000010011001101011",
						 "001001000010010111110110",
						 "001001000010010110000001",
						 "001001000010010100001100",
						 "001001000010010010010111",
						 "001001000010010000100010",
						 "001001000010001110101101",
						 "001001000010001100111000",
						 "001001000010001011000011",
						 "001001000010001001001110",
						 "001001000010000111011001",
						 "001001000010000101100100",
						 "001001000010000011101111",
						 "001001000010000001111010",
						 "001001000010011101010101",
						 "001001000010011011100000",
						 "001001000010011001101011",
						 "001001000010010111110110",
						 "001001000010010110000001",
						 "001001000010010100001100",
						 "001001000010010010010111",
						 "001001000010010000100010",
						 "001001000010001110101101",
						 "001001000010001100111000",
						 "001001000010001011000011",
						 "001001000010001001001110",
						 "001001000010000111011001",
						 "001001000010000101100100",
						 "001001000010000011101111",
						 "001001000010000001111010",
						 "001000111111111010010111",
						 "001000111111111000100010",
						 "001000111111110110101101",
						 "001000111111110100111000",
						 "001000111111110011000011",
						 "001000111111110001001110",
						 "001000111111101111011001",
						 "001000111111101101100100",
						 "001000111111101011101111",
						 "001000111111101001111010",
						 "001000111111101000000101",
						 "001000111111100110010000",
						 "001000111111100100011011",
						 "001000111111100010100110",
						 "001000111111100000110001",
						 "001000111111011110111100",
						 "001000111111111010100110",
						 "001000111111111000110000",
						 "001000111111110110111010",
						 "001000111111110101000100",
						 "001000111111110011001110",
						 "001000111111110001011000",
						 "001000111111101111100010",
						 "001000111111101101101100",
						 "001000111111101011110110",
						 "001000111111101010000000",
						 "001000111111101000001010",
						 "001000111111100110010100",
						 "001000111111100100011110",
						 "001000111111100010101000",
						 "001000111111100000110010",
						 "001000111111011110111100",
						 "001000111111111010100110",
						 "001000111111111000110000",
						 "001000111111110110111010",
						 "001000111111110101000100",
						 "001000111111110011001110",
						 "001000111111110001011000",
						 "001000111111101111100010",
						 "001000111111101101101100",
						 "001000111111101011110110",
						 "001000111111101010000000",
						 "001000111111101000001010",
						 "001000111111100110010100",
						 "001000111111100100011110",
						 "001000111111100010101000",
						 "001000111111100000110010",
						 "001000111111011110111100",
						 "001000111111111010100110",
						 "001000111111111000110000",
						 "001000111111110110111010",
						 "001000111111110101000100",
						 "001000111111110011001110",
						 "001000111111110001011000",
						 "001000111111101111100010",
						 "001000111111101101101100",
						 "001000111111101011110110",
						 "001000111111101010000000",
						 "001000111111101000001010",
						 "001000111111100110010100",
						 "001000111111100100011110",
						 "001000111111100010101000",
						 "001000111111100000110010",
						 "001000111111011110111100",
						 "001000111111111010110101",
						 "001000111111111000111110",
						 "001000111111110111000111",
						 "001000111111110101010000",
						 "001000111111110011011001",
						 "001000111111110001100010",
						 "001000111111101111101011",
						 "001000111111101101110100",
						 "001000111111101011111101",
						 "001000111111101010000110",
						 "001000111111101000001111",
						 "001000111111100110011000",
						 "001000111111100100100001",
						 "001000111111100010101010",
						 "001000111111100000110011",
						 "001000111111011110111100",
						 "001000111101010111110111",
						 "001000111101010110000000",
						 "001000111101010100001001",
						 "001000111101010010010010",
						 "001000111101010000011011",
						 "001000111101001110100100",
						 "001000111101001100101101",
						 "001000111101001010110110",
						 "001000111101001000111111",
						 "001000111101000111001000",
						 "001000111101000101010001",
						 "001000111101000011011010",
						 "001000111101000001100011",
						 "001000111100111111101100",
						 "001000111100111101110101",
						 "001000111100111011111110",
						 "001000111101010111110111",
						 "001000111101010110000000",
						 "001000111101010100001001",
						 "001000111101010010010010",
						 "001000111101010000011011",
						 "001000111101001110100100",
						 "001000111101001100101101",
						 "001000111101001010110110",
						 "001000111101001000111111",
						 "001000111101000111001000",
						 "001000111101000101010001",
						 "001000111101000011011010",
						 "001000111101000001100011",
						 "001000111100111111101100",
						 "001000111100111101110101",
						 "001000111100111011111110",
						 "001000111101011000000110",
						 "001000111101010110001110",
						 "001000111101010100010110",
						 "001000111101010010011110",
						 "001000111101010000100110",
						 "001000111101001110101110",
						 "001000111101001100110110",
						 "001000111101001010111110",
						 "001000111101001001000110",
						 "001000111101000111001110",
						 "001000111101000101010110",
						 "001000111101000011011110",
						 "001000111101000001100110",
						 "001000111100111111101110",
						 "001000111100111101110110",
						 "001000111100111011111110",
						 "001000111101011000000110",
						 "001000111101010110001110",
						 "001000111101010100010110",
						 "001000111101010010011110",
						 "001000111101010000100110",
						 "001000111101001110101110",
						 "001000111101001100110110",
						 "001000111101001010111110",
						 "001000111101001001000110",
						 "001000111101000111001110",
						 "001000111101000101010110",
						 "001000111101000011011110",
						 "001000111101000001100110",
						 "001000111100111111101110",
						 "001000111100111101110110",
						 "001000111100111011111110",
						 "001000111101011000000110",
						 "001000111101010110001110",
						 "001000111101010100010110",
						 "001000111101010010011110",
						 "001000111101010000100110",
						 "001000111101001110101110",
						 "001000111101001100110110",
						 "001000111101001010111110",
						 "001000111101001001000110",
						 "001000111101000111001110",
						 "001000111101000101010110",
						 "001000111101000011011110",
						 "001000111101000001100110",
						 "001000111100111111101110",
						 "001000111100111101110110",
						 "001000111100111011111110",
						 "001000111101011000010101",
						 "001000111101010110011100",
						 "001000111101010100100011",
						 "001000111101010010101010",
						 "001000111101010000110001",
						 "001000111101001110111000",
						 "001000111101001100111111",
						 "001000111101001011000110",
						 "001000111101001001001101",
						 "001000111101000111010100",
						 "001000111101000101011011",
						 "001000111101000011100010",
						 "001000111101000001101001",
						 "001000111100111111110000",
						 "001000111100111101110111",
						 "001000111100111011111110",
						 "001000111010110101010111",
						 "001000111010110011011110",
						 "001000111010110001100101",
						 "001000111010101111101100",
						 "001000111010101101110011",
						 "001000111010101011111010",
						 "001000111010101010000001",
						 "001000111010101000001000",
						 "001000111010100110001111",
						 "001000111010100100010110",
						 "001000111010100010011101",
						 "001000111010100000100100",
						 "001000111010011110101011",
						 "001000111010011100110010",
						 "001000111010011010111001",
						 "001000111010011001000000",
						 "001000111010110101010111",
						 "001000111010110011011110",
						 "001000111010110001100101",
						 "001000111010101111101100",
						 "001000111010101101110011",
						 "001000111010101011111010",
						 "001000111010101010000001",
						 "001000111010101000001000",
						 "001000111010100110001111",
						 "001000111010100100010110",
						 "001000111010100010011101",
						 "001000111010100000100100",
						 "001000111010011110101011",
						 "001000111010011100110010",
						 "001000111010011010111001",
						 "001000111010011001000000",
						 "001000111010110101100110",
						 "001000111010110011101100",
						 "001000111010110001110010",
						 "001000111010101111111000",
						 "001000111010101101111110",
						 "001000111010101100000100",
						 "001000111010101010001010",
						 "001000111010101000010000",
						 "001000111010100110010110",
						 "001000111010100100011100",
						 "001000111010100010100010",
						 "001000111010100000101000",
						 "001000111010011110101110",
						 "001000111010011100110100",
						 "001000111010011010111010",
						 "001000111010011001000000",
						 "001000111010110101100110",
						 "001000111010110011101100",
						 "001000111010110001110010",
						 "001000111010101111111000",
						 "001000111010101101111110",
						 "001000111010101100000100",
						 "001000111010101010001010",
						 "001000111010101000010000",
						 "001000111010100110010110",
						 "001000111010100100011100",
						 "001000111010100010100010",
						 "001000111010100000101000",
						 "001000111010011110101110",
						 "001000111010011100110100",
						 "001000111010011010111010",
						 "001000111010011001000000",
						 "001000111010110101100110",
						 "001000111010110011101100",
						 "001000111010110001110010",
						 "001000111010101111111000",
						 "001000111010101101111110",
						 "001000111010101100000100",
						 "001000111010101010001010",
						 "001000111010101000010000",
						 "001000111010100110010110",
						 "001000111010100100011100",
						 "001000111010100010100010",
						 "001000111010100000101000",
						 "001000111010011110101110",
						 "001000111010011100110100",
						 "001000111010011010111010",
						 "001000111010011001000000",
						 "001000111000010010110111",
						 "001000111000010000111100",
						 "001000111000001111000001",
						 "001000111000001101000110",
						 "001000111000001011001011",
						 "001000111000001001010000",
						 "001000111000000111010101",
						 "001000111000000101011010",
						 "001000111000000011011111",
						 "001000111000000001100100",
						 "001000110111111111101001",
						 "001000110111111101101110",
						 "001000110111111011110011",
						 "001000110111111001111000",
						 "001000110111110111111101",
						 "001000110111110110000010",
						 "001000111000010010110111",
						 "001000111000010000111100",
						 "001000111000001111000001",
						 "001000111000001101000110",
						 "001000111000001011001011",
						 "001000111000001001010000",
						 "001000111000000111010101",
						 "001000111000000101011010",
						 "001000111000000011011111",
						 "001000111000000001100100",
						 "001000110111111111101001",
						 "001000110111111101101110",
						 "001000110111111011110011",
						 "001000110111111001111000",
						 "001000110111110111111101",
						 "001000110111110110000010",
						 "001000111000010010110111",
						 "001000111000010000111100",
						 "001000111000001111000001",
						 "001000111000001101000110",
						 "001000111000001011001011",
						 "001000111000001001010000",
						 "001000111000000111010101",
						 "001000111000000101011010",
						 "001000111000000011011111",
						 "001000111000000001100100",
						 "001000110111111111101001",
						 "001000110111111101101110",
						 "001000110111111011110011",
						 "001000110111111001111000",
						 "001000110111110111111101",
						 "001000110111110110000010",
						 "001000111000010011000110",
						 "001000111000010001001010",
						 "001000111000001111001110",
						 "001000111000001101010010",
						 "001000111000001011010110",
						 "001000111000001001011010",
						 "001000111000000111011110",
						 "001000111000000101100010",
						 "001000111000000011100110",
						 "001000111000000001101010",
						 "001000110111111111101110",
						 "001000110111111101110010",
						 "001000110111111011110110",
						 "001000110111111001111010",
						 "001000110111110111111110",
						 "001000110111110110000010",
						 "001000111000010011000110",
						 "001000111000010001001010",
						 "001000111000001111001110",
						 "001000111000001101010010",
						 "001000111000001011010110",
						 "001000111000001001011010",
						 "001000111000000111011110",
						 "001000111000000101100010",
						 "001000111000000011100110",
						 "001000111000000001101010",
						 "001000110111111111101110",
						 "001000110111111101110010",
						 "001000110111111011110110",
						 "001000110111111001111010",
						 "001000110111110111111110",
						 "001000110111110110000010",
						 "001000110101110000001000",
						 "001000110101101110001100",
						 "001000110101101100010000",
						 "001000110101101010010100",
						 "001000110101101000011000",
						 "001000110101100110011100",
						 "001000110101100100100000",
						 "001000110101100010100100",
						 "001000110101100000101000",
						 "001000110101011110101100",
						 "001000110101011100110000",
						 "001000110101011010110100",
						 "001000110101011000111000",
						 "001000110101010110111100",
						 "001000110101010101000000",
						 "001000110101010011000100",
						 "001000110101110000010111",
						 "001000110101101110011010",
						 "001000110101101100011101",
						 "001000110101101010100000",
						 "001000110101101000100011",
						 "001000110101100110100110",
						 "001000110101100100101001",
						 "001000110101100010101100",
						 "001000110101100000101111",
						 "001000110101011110110010",
						 "001000110101011100110101",
						 "001000110101011010111000",
						 "001000110101011000111011",
						 "001000110101010110111110",
						 "001000110101010101000001",
						 "001000110101010011000100",
						 "001000110101110000010111",
						 "001000110101101110011010",
						 "001000110101101100011101",
						 "001000110101101010100000",
						 "001000110101101000100011",
						 "001000110101100110100110",
						 "001000110101100100101001",
						 "001000110101100010101100",
						 "001000110101100000101111",
						 "001000110101011110110010",
						 "001000110101011100110101",
						 "001000110101011010111000",
						 "001000110101011000111011",
						 "001000110101010110111110",
						 "001000110101010101000001",
						 "001000110101010011000100",
						 "001000110101110000100110",
						 "001000110101101110101000",
						 "001000110101101100101010",
						 "001000110101101010101100",
						 "001000110101101000101110",
						 "001000110101100110110000",
						 "001000110101100100110010",
						 "001000110101100010110100",
						 "001000110101100000110110",
						 "001000110101011110111000",
						 "001000110101011100111010",
						 "001000110101011010111100",
						 "001000110101011000111110",
						 "001000110101010111000000",
						 "001000110101010101000010",
						 "001000110101010011000100",
						 "001000110101110000100110",
						 "001000110101101110101000",
						 "001000110101101100101010",
						 "001000110101101010101100",
						 "001000110101101000101110",
						 "001000110101100110110000",
						 "001000110101100100110010",
						 "001000110101100010110100",
						 "001000110101100000110110",
						 "001000110101011110111000",
						 "001000110101011100111010",
						 "001000110101011010111100",
						 "001000110101011000111110",
						 "001000110101010111000000",
						 "001000110101010101000010",
						 "001000110101010011000100",
						 "001000110011001101101000",
						 "001000110011001011101010",
						 "001000110011001001101100",
						 "001000110011000111101110",
						 "001000110011000101110000",
						 "001000110011000011110010",
						 "001000110011000001110100",
						 "001000110010111111110110",
						 "001000110010111101111000",
						 "001000110010111011111010",
						 "001000110010111001111100",
						 "001000110010110111111110",
						 "001000110010110110000000",
						 "001000110010110100000010",
						 "001000110010110010000100",
						 "001000110010110000000110",
						 "001000110011001101110111",
						 "001000110011001011111000",
						 "001000110011001001111001",
						 "001000110011000111111010",
						 "001000110011000101111011",
						 "001000110011000011111100",
						 "001000110011000001111101",
						 "001000110010111111111110",
						 "001000110010111101111111",
						 "001000110010111100000000",
						 "001000110010111010000001",
						 "001000110010111000000010",
						 "001000110010110110000011",
						 "001000110010110100000100",
						 "001000110010110010000101",
						 "001000110010110000000110",
						 "001000110011001101110111",
						 "001000110011001011111000",
						 "001000110011001001111001",
						 "001000110011000111111010",
						 "001000110011000101111011",
						 "001000110011000011111100",
						 "001000110011000001111101",
						 "001000110010111111111110",
						 "001000110010111101111111",
						 "001000110010111100000000",
						 "001000110010111010000001",
						 "001000110010111000000010",
						 "001000110010110110000011",
						 "001000110010110100000100",
						 "001000110010110010000101",
						 "001000110010110000000110",
						 "001000110011001101110111",
						 "001000110011001011111000",
						 "001000110011001001111001",
						 "001000110011000111111010",
						 "001000110011000101111011",
						 "001000110011000011111100",
						 "001000110011000001111101",
						 "001000110010111111111110",
						 "001000110010111101111111",
						 "001000110010111100000000",
						 "001000110010111010000001",
						 "001000110010111000000010",
						 "001000110010110110000011",
						 "001000110010110100000100",
						 "001000110010110010000101",
						 "001000110010110000000110",
						 "001000110011001110000110",
						 "001000110011001100000110",
						 "001000110011001010000110",
						 "001000110011001000000110",
						 "001000110011000110000110",
						 "001000110011000100000110",
						 "001000110011000010000110",
						 "001000110011000000000110",
						 "001000110010111110000110",
						 "001000110010111100000110",
						 "001000110010111010000110",
						 "001000110010111000000110",
						 "001000110010110110000110",
						 "001000110010110100000110",
						 "001000110010110010000110",
						 "001000110010110000000110",
						 "001000110011001110000110",
						 "001000110011001100000110",
						 "001000110011001010000110",
						 "001000110011001000000110",
						 "001000110011000110000110",
						 "001000110011000100000110",
						 "001000110011000010000110",
						 "001000110011000000000110",
						 "001000110010111110000110",
						 "001000110010111100000110",
						 "001000110010111010000110",
						 "001000110010111000000110",
						 "001000110010110110000110",
						 "001000110010110100000110",
						 "001000110010110010000110",
						 "001000110010110000000110",
						 "001000110000101011001000",
						 "001000110000101001001000",
						 "001000110000100111001000",
						 "001000110000100101001000",
						 "001000110000100011001000",
						 "001000110000100001001000",
						 "001000110000011111001000",
						 "001000110000011101001000",
						 "001000110000011011001000",
						 "001000110000011001001000",
						 "001000110000010111001000",
						 "001000110000010101001000",
						 "001000110000010011001000",
						 "001000110000010001001000",
						 "001000110000001111001000",
						 "001000110000001101001000",
						 "001000110000101011010111",
						 "001000110000101001010110",
						 "001000110000100111010101",
						 "001000110000100101010100",
						 "001000110000100011010011",
						 "001000110000100001010010",
						 "001000110000011111010001",
						 "001000110000011101010000",
						 "001000110000011011001111",
						 "001000110000011001001110",
						 "001000110000010111001101",
						 "001000110000010101001100",
						 "001000110000010011001011",
						 "001000110000010001001010",
						 "001000110000001111001001",
						 "001000110000001101001000",
						 "001000110000101011010111",
						 "001000110000101001010110",
						 "001000110000100111010101",
						 "001000110000100101010100",
						 "001000110000100011010011",
						 "001000110000100001010010",
						 "001000110000011111010001",
						 "001000110000011101010000",
						 "001000110000011011001111",
						 "001000110000011001001110",
						 "001000110000010111001101",
						 "001000110000010101001100",
						 "001000110000010011001011",
						 "001000110000010001001010",
						 "001000110000001111001001",
						 "001000110000001101001000",
						 "001000110000101011010111",
						 "001000110000101001010110",
						 "001000110000100111010101",
						 "001000110000100101010100",
						 "001000110000100011010011",
						 "001000110000100001010010",
						 "001000110000011111010001",
						 "001000110000011101010000",
						 "001000110000011011001111",
						 "001000110000011001001110",
						 "001000110000010111001101",
						 "001000110000010101001100",
						 "001000110000010011001011",
						 "001000110000010001001010",
						 "001000110000001111001001",
						 "001000110000001101001000",
						 "001000110000101011100110",
						 "001000110000101001100100",
						 "001000110000100111100010",
						 "001000110000100101100000",
						 "001000110000100011011110",
						 "001000110000100001011100",
						 "001000110000011111011010",
						 "001000110000011101011000",
						 "001000110000011011010110",
						 "001000110000011001010100",
						 "001000110000010111010010",
						 "001000110000010101010000",
						 "001000110000010011001110",
						 "001000110000010001001100",
						 "001000110000001111001010",
						 "001000110000001101001000",
						 "001000101110001000101000",
						 "001000101110000110100110",
						 "001000101110000100100100",
						 "001000101110000010100010",
						 "001000101110000000100000",
						 "001000101101111110011110",
						 "001000101101111100011100",
						 "001000101101111010011010",
						 "001000101101111000011000",
						 "001000101101110110010110",
						 "001000101101110100010100",
						 "001000101101110010010010",
						 "001000101101110000010000",
						 "001000101101101110001110",
						 "001000101101101100001100",
						 "001000101101101010001010",
						 "001000101110001000101000",
						 "001000101110000110100110",
						 "001000101110000100100100",
						 "001000101110000010100010",
						 "001000101110000000100000",
						 "001000101101111110011110",
						 "001000101101111100011100",
						 "001000101101111010011010",
						 "001000101101111000011000",
						 "001000101101110110010110",
						 "001000101101110100010100",
						 "001000101101110010010010",
						 "001000101101110000010000",
						 "001000101101101110001110",
						 "001000101101101100001100",
						 "001000101101101010001010",
						 "001000101110001000110111",
						 "001000101110000110110100",
						 "001000101110000100110001",
						 "001000101110000010101110",
						 "001000101110000000101011",
						 "001000101101111110101000",
						 "001000101101111100100101",
						 "001000101101111010100010",
						 "001000101101111000011111",
						 "001000101101110110011100",
						 "001000101101110100011001",
						 "001000101101110010010110",
						 "001000101101110000010011",
						 "001000101101101110010000",
						 "001000101101101100001101",
						 "001000101101101010001010",
						 "001000101110001000110111",
						 "001000101110000110110100",
						 "001000101110000100110001",
						 "001000101110000010101110",
						 "001000101110000000101011",
						 "001000101101111110101000",
						 "001000101101111100100101",
						 "001000101101111010100010",
						 "001000101101111000011111",
						 "001000101101110110011100",
						 "001000101101110100011001",
						 "001000101101110010010110",
						 "001000101101110000010011",
						 "001000101101101110010000",
						 "001000101101101100001101",
						 "001000101101101010001010",
						 "001000101110001000110111",
						 "001000101110000110110100",
						 "001000101110000100110001",
						 "001000101110000010101110",
						 "001000101110000000101011",
						 "001000101101111110101000",
						 "001000101101111100100101",
						 "001000101101111010100010",
						 "001000101101111000011111",
						 "001000101101110110011100",
						 "001000101101110100011001",
						 "001000101101110010010110",
						 "001000101101110000010011",
						 "001000101101101110010000",
						 "001000101101101100001101",
						 "001000101101101010001010",
						 "001000101011100110001000",
						 "001000101011100100000100",
						 "001000101011100010000000",
						 "001000101011011111111100",
						 "001000101011011101111000",
						 "001000101011011011110100",
						 "001000101011011001110000",
						 "001000101011010111101100",
						 "001000101011010101101000",
						 "001000101011010011100100",
						 "001000101011010001100000",
						 "001000101011001111011100",
						 "001000101011001101011000",
						 "001000101011001011010100",
						 "001000101011001001010000",
						 "001000101011000111001100",
						 "001000101011100110001000",
						 "001000101011100100000100",
						 "001000101011100010000000",
						 "001000101011011111111100",
						 "001000101011011101111000",
						 "001000101011011011110100",
						 "001000101011011001110000",
						 "001000101011010111101100",
						 "001000101011010101101000",
						 "001000101011010011100100",
						 "001000101011010001100000",
						 "001000101011001111011100",
						 "001000101011001101011000",
						 "001000101011001011010100",
						 "001000101011001001010000",
						 "001000101011000111001100",
						 "001000101011100110001000",
						 "001000101011100100000100",
						 "001000101011100010000000",
						 "001000101011011111111100",
						 "001000101011011101111000",
						 "001000101011011011110100",
						 "001000101011011001110000",
						 "001000101011010111101100",
						 "001000101011010101101000",
						 "001000101011010011100100",
						 "001000101011010001100000",
						 "001000101011001111011100",
						 "001000101011001101011000",
						 "001000101011001011010100",
						 "001000101011001001010000",
						 "001000101011000111001100",
						 "001000101011100110010111",
						 "001000101011100100010010",
						 "001000101011100010001101",
						 "001000101011100000001000",
						 "001000101011011110000011",
						 "001000101011011011111110",
						 "001000101011011001111001",
						 "001000101011010111110100",
						 "001000101011010101101111",
						 "001000101011010011101010",
						 "001000101011010001100101",
						 "001000101011001111100000",
						 "001000101011001101011011",
						 "001000101011001011010110",
						 "001000101011001001010001",
						 "001000101011000111001100",
						 "001000101011100110010111",
						 "001000101011100100010010",
						 "001000101011100010001101",
						 "001000101011100000001000",
						 "001000101011011110000011",
						 "001000101011011011111110",
						 "001000101011011001111001",
						 "001000101011010111110100",
						 "001000101011010101101111",
						 "001000101011010011101010",
						 "001000101011010001100101",
						 "001000101011001111100000",
						 "001000101011001101011011",
						 "001000101011001011010110",
						 "001000101011001001010001",
						 "001000101011000111001100",
						 "001000101001000011011001",
						 "001000101001000001010100",
						 "001000101000111111001111",
						 "001000101000111101001010",
						 "001000101000111011000101",
						 "001000101000111001000000",
						 "001000101000110110111011",
						 "001000101000110100110110",
						 "001000101000110010110001",
						 "001000101000110000101100",
						 "001000101000101110100111",
						 "001000101000101100100010",
						 "001000101000101010011101",
						 "001000101000101000011000",
						 "001000101000100110010011",
						 "001000101000100100001110",
						 "001000101001000011101000",
						 "001000101001000001100010",
						 "001000101000111111011100",
						 "001000101000111101010110",
						 "001000101000111011010000",
						 "001000101000111001001010",
						 "001000101000110111000100",
						 "001000101000110100111110",
						 "001000101000110010111000",
						 "001000101000110000110010",
						 "001000101000101110101100",
						 "001000101000101100100110",
						 "001000101000101010100000",
						 "001000101000101000011010",
						 "001000101000100110010100",
						 "001000101000100100001110",
						 "001000101001000011101000",
						 "001000101001000001100010",
						 "001000101000111111011100",
						 "001000101000111101010110",
						 "001000101000111011010000",
						 "001000101000111001001010",
						 "001000101000110111000100",
						 "001000101000110100111110",
						 "001000101000110010111000",
						 "001000101000110000110010",
						 "001000101000101110101100",
						 "001000101000101100100110",
						 "001000101000101010100000",
						 "001000101000101000011010",
						 "001000101000100110010100",
						 "001000101000100100001110",
						 "001000101001000011101000",
						 "001000101001000001100010",
						 "001000101000111111011100",
						 "001000101000111101010110",
						 "001000101000111011010000",
						 "001000101000111001001010",
						 "001000101000110111000100",
						 "001000101000110100111110",
						 "001000101000110010111000",
						 "001000101000110000110010",
						 "001000101000101110101100",
						 "001000101000101100100110",
						 "001000101000101010100000",
						 "001000101000101000011010",
						 "001000101000100110010100",
						 "001000101000100100001110",
						 "001000100110100000111001",
						 "001000100110011110110010",
						 "001000100110011100101011",
						 "001000100110011010100100",
						 "001000100110011000011101",
						 "001000100110010110010110",
						 "001000100110010100001111",
						 "001000100110010010001000",
						 "001000100110010000000001",
						 "001000100110001101111010",
						 "001000100110001011110011",
						 "001000100110001001101100",
						 "001000100110000111100101",
						 "001000100110000101011110",
						 "001000100110000011010111",
						 "001000100110000001010000",
						 "001000100110100000111001",
						 "001000100110011110110010",
						 "001000100110011100101011",
						 "001000100110011010100100",
						 "001000100110011000011101",
						 "001000100110010110010110",
						 "001000100110010100001111",
						 "001000100110010010001000",
						 "001000100110010000000001",
						 "001000100110001101111010",
						 "001000100110001011110011",
						 "001000100110001001101100",
						 "001000100110000111100101",
						 "001000100110000101011110",
						 "001000100110000011010111",
						 "001000100110000001010000",
						 "001000100110100000111001",
						 "001000100110011110110010",
						 "001000100110011100101011",
						 "001000100110011010100100",
						 "001000100110011000011101",
						 "001000100110010110010110",
						 "001000100110010100001111",
						 "001000100110010010001000",
						 "001000100110010000000001",
						 "001000100110001101111010",
						 "001000100110001011110011",
						 "001000100110001001101100",
						 "001000100110000111100101",
						 "001000100110000101011110",
						 "001000100110000011010111",
						 "001000100110000001010000",
						 "001000100110100001001000",
						 "001000100110011111000000",
						 "001000100110011100111000",
						 "001000100110011010110000",
						 "001000100110011000101000",
						 "001000100110010110100000",
						 "001000100110010100011000",
						 "001000100110010010010000",
						 "001000100110010000001000",
						 "001000100110001110000000",
						 "001000100110001011111000",
						 "001000100110001001110000",
						 "001000100110000111101000",
						 "001000100110000101100000",
						 "001000100110000011011000",
						 "001000100110000001010000",
						 "001000100110100001001000",
						 "001000100110011111000000",
						 "001000100110011100111000",
						 "001000100110011010110000",
						 "001000100110011000101000",
						 "001000100110010110100000",
						 "001000100110010100011000",
						 "001000100110010010010000",
						 "001000100110010000001000",
						 "001000100110001110000000",
						 "001000100110001011111000",
						 "001000100110001001110000",
						 "001000100110000111101000",
						 "001000100110000101100000",
						 "001000100110000011011000",
						 "001000100110000001010000",
						 "001000100011111110001010",
						 "001000100011111100000010",
						 "001000100011111001111010",
						 "001000100011110111110010",
						 "001000100011110101101010",
						 "001000100011110011100010",
						 "001000100011110001011010",
						 "001000100011101111010010",
						 "001000100011101101001010",
						 "001000100011101011000010",
						 "001000100011101000111010",
						 "001000100011100110110010",
						 "001000100011100100101010",
						 "001000100011100010100010",
						 "001000100011100000011010",
						 "001000100011011110010010",
						 "001000100011111110011001",
						 "001000100011111100010000",
						 "001000100011111010000111",
						 "001000100011110111111110",
						 "001000100011110101110101",
						 "001000100011110011101100",
						 "001000100011110001100011",
						 "001000100011101111011010",
						 "001000100011101101010001",
						 "001000100011101011001000",
						 "001000100011101000111111",
						 "001000100011100110110110",
						 "001000100011100100101101",
						 "001000100011100010100100",
						 "001000100011100000011011",
						 "001000100011011110010010",
						 "001000100011111110011001",
						 "001000100011111100010000",
						 "001000100011111010000111",
						 "001000100011110111111110",
						 "001000100011110101110101",
						 "001000100011110011101100",
						 "001000100011110001100011",
						 "001000100011101111011010",
						 "001000100011101101010001",
						 "001000100011101011001000",
						 "001000100011101000111111",
						 "001000100011100110110110",
						 "001000100011100100101101",
						 "001000100011100010100100",
						 "001000100011100000011011",
						 "001000100011011110010010",
						 "001000100011111110011001",
						 "001000100011111100010000",
						 "001000100011111010000111",
						 "001000100011110111111110",
						 "001000100011110101110101",
						 "001000100011110011101100",
						 "001000100011110001100011",
						 "001000100011101111011010",
						 "001000100011101101010001",
						 "001000100011101011001000",
						 "001000100011101000111111",
						 "001000100011100110110110",
						 "001000100011100100101101",
						 "001000100011100010100100",
						 "001000100011100000011011",
						 "001000100011011110010010",
						 "001000100011111110101000",
						 "001000100011111100011110",
						 "001000100011111010010100",
						 "001000100011111000001010",
						 "001000100011110110000000",
						 "001000100011110011110110",
						 "001000100011110001101100",
						 "001000100011101111100010",
						 "001000100011101101011000",
						 "001000100011101011001110",
						 "001000100011101001000100",
						 "001000100011100110111010",
						 "001000100011100100110000",
						 "001000100011100010100110",
						 "001000100011100000011100",
						 "001000100011011110010010",
						 "001000100001011011101010",
						 "001000100001011001100000",
						 "001000100001010111010110",
						 "001000100001010101001100",
						 "001000100001010011000010",
						 "001000100001010000111000",
						 "001000100001001110101110",
						 "001000100001001100100100",
						 "001000100001001010011010",
						 "001000100001001000010000",
						 "001000100001000110000110",
						 "001000100001000011111100",
						 "001000100001000001110010",
						 "001000100000111111101000",
						 "001000100000111101011110",
						 "001000100000111011010100",
						 "001000100001011011101010",
						 "001000100001011001100000",
						 "001000100001010111010110",
						 "001000100001010101001100",
						 "001000100001010011000010",
						 "001000100001010000111000",
						 "001000100001001110101110",
						 "001000100001001100100100",
						 "001000100001001010011010",
						 "001000100001001000010000",
						 "001000100001000110000110",
						 "001000100001000011111100",
						 "001000100001000001110010",
						 "001000100000111111101000",
						 "001000100000111101011110",
						 "001000100000111011010100",
						 "001000100001011011111001",
						 "001000100001011001101110",
						 "001000100001010111100011",
						 "001000100001010101011000",
						 "001000100001010011001101",
						 "001000100001010001000010",
						 "001000100001001110110111",
						 "001000100001001100101100",
						 "001000100001001010100001",
						 "001000100001001000010110",
						 "001000100001000110001011",
						 "001000100001000100000000",
						 "001000100001000001110101",
						 "001000100000111111101010",
						 "001000100000111101011111",
						 "001000100000111011010100",
						 "001000100001011011111001",
						 "001000100001011001101110",
						 "001000100001010111100011",
						 "001000100001010101011000",
						 "001000100001010011001101",
						 "001000100001010001000010",
						 "001000100001001110110111",
						 "001000100001001100101100",
						 "001000100001001010100001",
						 "001000100001001000010110",
						 "001000100001000110001011",
						 "001000100001000100000000",
						 "001000100001000001110101",
						 "001000100000111111101010",
						 "001000100000111101011111",
						 "001000100000111011010100",
						 "001000100001011011111001",
						 "001000100001011001101110",
						 "001000100001010111100011",
						 "001000100001010101011000",
						 "001000100001010011001101",
						 "001000100001010001000010",
						 "001000100001001110110111",
						 "001000100001001100101100",
						 "001000100001001010100001",
						 "001000100001001000010110",
						 "001000100001000110001011",
						 "001000100001000100000000",
						 "001000100001000001110101",
						 "001000100000111111101010",
						 "001000100000111101011111",
						 "001000100000111011010100",
						 "001000011110111001001010",
						 "001000011110110110111110",
						 "001000011110110100110010",
						 "001000011110110010100110",
						 "001000011110110000011010",
						 "001000011110101110001110",
						 "001000011110101100000010",
						 "001000011110101001110110",
						 "001000011110100111101010",
						 "001000011110100101011110",
						 "001000011110100011010010",
						 "001000011110100001000110",
						 "001000011110011110111010",
						 "001000011110011100101110",
						 "001000011110011010100010",
						 "001000011110011000010110",
						 "001000011110111001001010",
						 "001000011110110110111110",
						 "001000011110110100110010",
						 "001000011110110010100110",
						 "001000011110110000011010",
						 "001000011110101110001110",
						 "001000011110101100000010",
						 "001000011110101001110110",
						 "001000011110100111101010",
						 "001000011110100101011110",
						 "001000011110100011010010",
						 "001000011110100001000110",
						 "001000011110011110111010",
						 "001000011110011100101110",
						 "001000011110011010100010",
						 "001000011110011000010110",
						 "001000011110111001001010",
						 "001000011110110110111110",
						 "001000011110110100110010",
						 "001000011110110010100110",
						 "001000011110110000011010",
						 "001000011110101110001110",
						 "001000011110101100000010",
						 "001000011110101001110110",
						 "001000011110100111101010",
						 "001000011110100101011110",
						 "001000011110100011010010",
						 "001000011110100001000110",
						 "001000011110011110111010",
						 "001000011110011100101110",
						 "001000011110011010100010",
						 "001000011110011000010110",
						 "001000011110111001011001",
						 "001000011110110111001100",
						 "001000011110110100111111",
						 "001000011110110010110010",
						 "001000011110110000100101",
						 "001000011110101110011000",
						 "001000011110101100001011",
						 "001000011110101001111110",
						 "001000011110100111110001",
						 "001000011110100101100100",
						 "001000011110100011010111",
						 "001000011110100001001010",
						 "001000011110011110111101",
						 "001000011110011100110000",
						 "001000011110011010100011",
						 "001000011110011000010110",
						 "001000011100010110011011",
						 "001000011100010100001110",
						 "001000011100010010000001",
						 "001000011100001111110100",
						 "001000011100001101100111",
						 "001000011100001011011010",
						 "001000011100001001001101",
						 "001000011100000111000000",
						 "001000011100000100110011",
						 "001000011100000010100110",
						 "001000011100000000011001",
						 "001000011011111110001100",
						 "001000011011111011111111",
						 "001000011011111001110010",
						 "001000011011110111100101",
						 "001000011011110101011000",
						 "001000011100010110011011",
						 "001000011100010100001110",
						 "001000011100010010000001",
						 "001000011100001111110100",
						 "001000011100001101100111",
						 "001000011100001011011010",
						 "001000011100001001001101",
						 "001000011100000111000000",
						 "001000011100000100110011",
						 "001000011100000010100110",
						 "001000011100000000011001",
						 "001000011011111110001100",
						 "001000011011111011111111",
						 "001000011011111001110010",
						 "001000011011110111100101",
						 "001000011011110101011000",
						 "001000011100010110101010",
						 "001000011100010100011100",
						 "001000011100010010001110",
						 "001000011100010000000000",
						 "001000011100001101110010",
						 "001000011100001011100100",
						 "001000011100001001010110",
						 "001000011100000111001000",
						 "001000011100000100111010",
						 "001000011100000010101100",
						 "001000011100000000011110",
						 "001000011011111110010000",
						 "001000011011111100000010",
						 "001000011011111001110100",
						 "001000011011110111100110",
						 "001000011011110101011000",
						 "001000011100010110101010",
						 "001000011100010100011100",
						 "001000011100010010001110",
						 "001000011100010000000000",
						 "001000011100001101110010",
						 "001000011100001011100100",
						 "001000011100001001010110",
						 "001000011100000111001000",
						 "001000011100000100111010",
						 "001000011100000010101100",
						 "001000011100000000011110",
						 "001000011011111110010000",
						 "001000011011111100000010",
						 "001000011011111001110100",
						 "001000011011110111100110",
						 "001000011011110101011000",
						 "001000011100010110101010",
						 "001000011100010100011100",
						 "001000011100010010001110",
						 "001000011100010000000000",
						 "001000011100001101110010",
						 "001000011100001011100100",
						 "001000011100001001010110",
						 "001000011100000111001000",
						 "001000011100000100111010",
						 "001000011100000010101100",
						 "001000011100000000011110",
						 "001000011011111110010000",
						 "001000011011111100000010",
						 "001000011011111001110100",
						 "001000011011110111100110",
						 "001000011011110101011000",
						 "001000011001110011101100",
						 "001000011001110001011110",
						 "001000011001101111010000",
						 "001000011001101101000010",
						 "001000011001101010110100",
						 "001000011001101000100110",
						 "001000011001100110011000",
						 "001000011001100100001010",
						 "001000011001100001111100",
						 "001000011001011111101110",
						 "001000011001011101100000",
						 "001000011001011011010010",
						 "001000011001011001000100",
						 "001000011001010110110110",
						 "001000011001010100101000",
						 "001000011001010010011010",
						 "001000011001110011111011",
						 "001000011001110001101100",
						 "001000011001101111011101",
						 "001000011001101101001110",
						 "001000011001101010111111",
						 "001000011001101000110000",
						 "001000011001100110100001",
						 "001000011001100100010010",
						 "001000011001100010000011",
						 "001000011001011111110100",
						 "001000011001011101100101",
						 "001000011001011011010110",
						 "001000011001011001000111",
						 "001000011001010110111000",
						 "001000011001010100101001",
						 "001000011001010010011010",
						 "001000011001110011111011",
						 "001000011001110001101100",
						 "001000011001101111011101",
						 "001000011001101101001110",
						 "001000011001101010111111",
						 "001000011001101000110000",
						 "001000011001100110100001",
						 "001000011001100100010010",
						 "001000011001100010000011",
						 "001000011001011111110100",
						 "001000011001011101100101",
						 "001000011001011011010110",
						 "001000011001011001000111",
						 "001000011001010110111000",
						 "001000011001010100101001",
						 "001000011001010010011010",
						 "001000011001110011111011",
						 "001000011001110001101100",
						 "001000011001101111011101",
						 "001000011001101101001110",
						 "001000011001101010111111",
						 "001000011001101000110000",
						 "001000011001100110100001",
						 "001000011001100100010010",
						 "001000011001100010000011",
						 "001000011001011111110100",
						 "001000011001011101100101",
						 "001000011001011011010110",
						 "001000011001011001000111",
						 "001000011001010110111000",
						 "001000011001010100101001",
						 "001000011001010010011010",
						 "001000010111010001001100",
						 "001000010111001110111100",
						 "001000010111001100101100",
						 "001000010111001010011100",
						 "001000010111001000001100",
						 "001000010111000101111100",
						 "001000010111000011101100",
						 "001000010111000001011100",
						 "001000010110111111001100",
						 "001000010110111100111100",
						 "001000010110111010101100",
						 "001000010110111000011100",
						 "001000010110110110001100",
						 "001000010110110011111100",
						 "001000010110110001101100",
						 "001000010110101111011100",
						 "001000010111010001001100",
						 "001000010111001110111100",
						 "001000010111001100101100",
						 "001000010111001010011100",
						 "001000010111001000001100",
						 "001000010111000101111100",
						 "001000010111000011101100",
						 "001000010111000001011100",
						 "001000010110111111001100",
						 "001000010110111100111100",
						 "001000010110111010101100",
						 "001000010110111000011100",
						 "001000010110110110001100",
						 "001000010110110011111100",
						 "001000010110110001101100",
						 "001000010110101111011100",
						 "001000010111010001001100",
						 "001000010111001110111100",
						 "001000010111001100101100",
						 "001000010111001010011100",
						 "001000010111001000001100",
						 "001000010111000101111100",
						 "001000010111000011101100",
						 "001000010111000001011100",
						 "001000010110111111001100",
						 "001000010110111100111100",
						 "001000010110111010101100",
						 "001000010110111000011100",
						 "001000010110110110001100",
						 "001000010110110011111100",
						 "001000010110110001101100",
						 "001000010110101111011100",
						 "001000010111010001011011",
						 "001000010111001111001010",
						 "001000010111001100111001",
						 "001000010111001010101000",
						 "001000010111001000010111",
						 "001000010111000110000110",
						 "001000010111000011110101",
						 "001000010111000001100100",
						 "001000010110111111010011",
						 "001000010110111101000010",
						 "001000010110111010110001",
						 "001000010110111000100000",
						 "001000010110110110001111",
						 "001000010110110011111110",
						 "001000010110110001101101",
						 "001000010110101111011100",
						 "001000010111010001011011",
						 "001000010111001111001010",
						 "001000010111001100111001",
						 "001000010111001010101000",
						 "001000010111001000010111",
						 "001000010111000110000110",
						 "001000010111000011110101",
						 "001000010111000001100100",
						 "001000010110111111010011",
						 "001000010110111101000010",
						 "001000010110111010110001",
						 "001000010110111000100000",
						 "001000010110110110001111",
						 "001000010110110011111110",
						 "001000010110110001101101",
						 "001000010110101111011100",
						 "001000010100101110011101",
						 "001000010100101100001100",
						 "001000010100101001111011",
						 "001000010100100111101010",
						 "001000010100100101011001",
						 "001000010100100011001000",
						 "001000010100100000110111",
						 "001000010100011110100110",
						 "001000010100011100010101",
						 "001000010100011010000100",
						 "001000010100010111110011",
						 "001000010100010101100010",
						 "001000010100010011010001",
						 "001000010100010001000000",
						 "001000010100001110101111",
						 "001000010100001100011110",
						 "001000010100101110101100",
						 "001000010100101100011010",
						 "001000010100101010001000",
						 "001000010100100111110110",
						 "001000010100100101100100",
						 "001000010100100011010010",
						 "001000010100100001000000",
						 "001000010100011110101110",
						 "001000010100011100011100",
						 "001000010100011010001010",
						 "001000010100010111111000",
						 "001000010100010101100110",
						 "001000010100010011010100",
						 "001000010100010001000010",
						 "001000010100001110110000",
						 "001000010100001100011110",
						 "001000010100101110101100",
						 "001000010100101100011010",
						 "001000010100101010001000",
						 "001000010100100111110110",
						 "001000010100100101100100",
						 "001000010100100011010010",
						 "001000010100100001000000",
						 "001000010100011110101110",
						 "001000010100011100011100",
						 "001000010100011010001010",
						 "001000010100010111111000",
						 "001000010100010101100110",
						 "001000010100010011010100",
						 "001000010100010001000010",
						 "001000010100001110110000",
						 "001000010100001100011110",
						 "001000010100101110101100",
						 "001000010100101100011010",
						 "001000010100101010001000",
						 "001000010100100111110110",
						 "001000010100100101100100",
						 "001000010100100011010010",
						 "001000010100100001000000",
						 "001000010100011110101110",
						 "001000010100011100011100",
						 "001000010100011010001010",
						 "001000010100010111111000",
						 "001000010100010101100110",
						 "001000010100010011010100",
						 "001000010100010001000010",
						 "001000010100001110110000",
						 "001000010100001100011110",
						 "001000010010001011111101",
						 "001000010010001001101010",
						 "001000010010000111010111",
						 "001000010010000101000100",
						 "001000010010000010110001",
						 "001000010010000000011110",
						 "001000010001111110001011",
						 "001000010001111011111000",
						 "001000010001111001100101",
						 "001000010001110111010010",
						 "001000010001110100111111",
						 "001000010001110010101100",
						 "001000010001110000011001",
						 "001000010001101110000110",
						 "001000010001101011110011",
						 "001000010001101001100000",
						 "001000010010001011111101",
						 "001000010010001001101010",
						 "001000010010000111010111",
						 "001000010010000101000100",
						 "001000010010000010110001",
						 "001000010010000000011110",
						 "001000010001111110001011",
						 "001000010001111011111000",
						 "001000010001111001100101",
						 "001000010001110111010010",
						 "001000010001110100111111",
						 "001000010001110010101100",
						 "001000010001110000011001",
						 "001000010001101110000110",
						 "001000010001101011110011",
						 "001000010001101001100000",
						 "001000010010001011111101",
						 "001000010010001001101010",
						 "001000010010000111010111",
						 "001000010010000101000100",
						 "001000010010000010110001",
						 "001000010010000000011110",
						 "001000010001111110001011",
						 "001000010001111011111000",
						 "001000010001111001100101",
						 "001000010001110111010010",
						 "001000010001110100111111",
						 "001000010001110010101100",
						 "001000010001110000011001",
						 "001000010001101110000110",
						 "001000010001101011110011",
						 "001000010001101001100000",
						 "001000010010001100001100",
						 "001000010010001001111000",
						 "001000010010000111100100",
						 "001000010010000101010000",
						 "001000010010000010111100",
						 "001000010010000000101000",
						 "001000010001111110010100",
						 "001000010001111100000000",
						 "001000010001111001101100",
						 "001000010001110111011000",
						 "001000010001110101000100",
						 "001000010001110010110000",
						 "001000010001110000011100",
						 "001000010001101110001000",
						 "001000010001101011110100",
						 "001000010001101001100000",
						 "001000010010001100001100",
						 "001000010010001001111000",
						 "001000010010000111100100",
						 "001000010010000101010000",
						 "001000010010000010111100",
						 "001000010010000000101000",
						 "001000010001111110010100",
						 "001000010001111100000000",
						 "001000010001111001101100",
						 "001000010001110111011000",
						 "001000010001110101000100",
						 "001000010001110010110000",
						 "001000010001110000011100",
						 "001000010001101110001000",
						 "001000010001101011110100",
						 "001000010001101001100000",
						 "001000001111101001001110",
						 "001000001111100110111010",
						 "001000001111100100100110",
						 "001000001111100010010010",
						 "001000001111011111111110",
						 "001000001111011101101010",
						 "001000001111011011010110",
						 "001000001111011001000010",
						 "001000001111010110101110",
						 "001000001111010100011010",
						 "001000001111010010000110",
						 "001000001111001111110010",
						 "001000001111001101011110",
						 "001000001111001011001010",
						 "001000001111001000110110",
						 "001000001111000110100010",
						 "001000001111101001011101",
						 "001000001111100111001000",
						 "001000001111100100110011",
						 "001000001111100010011110",
						 "001000001111100000001001",
						 "001000001111011101110100",
						 "001000001111011011011111",
						 "001000001111011001001010",
						 "001000001111010110110101",
						 "001000001111010100100000",
						 "001000001111010010001011",
						 "001000001111001111110110",
						 "001000001111001101100001",
						 "001000001111001011001100",
						 "001000001111001000110111",
						 "001000001111000110100010",
						 "001000001111101001011101",
						 "001000001111100111001000",
						 "001000001111100100110011",
						 "001000001111100010011110",
						 "001000001111100000001001",
						 "001000001111011101110100",
						 "001000001111011011011111",
						 "001000001111011001001010",
						 "001000001111010110110101",
						 "001000001111010100100000",
						 "001000001111010010001011",
						 "001000001111001111110110",
						 "001000001111001101100001",
						 "001000001111001011001100",
						 "001000001111001000110111",
						 "001000001111000110100010",
						 "001000001111101001011101",
						 "001000001111100111001000",
						 "001000001111100100110011",
						 "001000001111100010011110",
						 "001000001111100000001001",
						 "001000001111011101110100",
						 "001000001111011011011111",
						 "001000001111011001001010",
						 "001000001111010110110101",
						 "001000001111010100100000",
						 "001000001111010010001011",
						 "001000001111001111110110",
						 "001000001111001101100001",
						 "001000001111001011001100",
						 "001000001111001000110111",
						 "001000001111000110100010",
						 "001000001101000110101110",
						 "001000001101000100011000",
						 "001000001101000010000010",
						 "001000001100111111101100",
						 "001000001100111101010110",
						 "001000001100111011000000",
						 "001000001100111000101010",
						 "001000001100110110010100",
						 "001000001100110011111110",
						 "001000001100110001101000",
						 "001000001100101111010010",
						 "001000001100101100111100",
						 "001000001100101010100110",
						 "001000001100101000010000",
						 "001000001100100101111010",
						 "001000001100100011100100",
						 "001000001101000110101110",
						 "001000001101000100011000",
						 "001000001101000010000010",
						 "001000001100111111101100",
						 "001000001100111101010110",
						 "001000001100111011000000",
						 "001000001100111000101010",
						 "001000001100110110010100",
						 "001000001100110011111110",
						 "001000001100110001101000",
						 "001000001100101111010010",
						 "001000001100101100111100",
						 "001000001100101010100110",
						 "001000001100101000010000",
						 "001000001100100101111010",
						 "001000001100100011100100",
						 "001000001101000110101110",
						 "001000001101000100011000",
						 "001000001101000010000010",
						 "001000001100111111101100",
						 "001000001100111101010110",
						 "001000001100111011000000",
						 "001000001100111000101010",
						 "001000001100110110010100",
						 "001000001100110011111110",
						 "001000001100110001101000",
						 "001000001100101111010010",
						 "001000001100101100111100",
						 "001000001100101010100110",
						 "001000001100101000010000",
						 "001000001100100101111010",
						 "001000001100100011100100",
						 "001000001101000110101110",
						 "001000001101000100011000",
						 "001000001101000010000010",
						 "001000001100111111101100",
						 "001000001100111101010110",
						 "001000001100111011000000",
						 "001000001100111000101010",
						 "001000001100110110010100",
						 "001000001100110011111110",
						 "001000001100110001101000",
						 "001000001100101111010010",
						 "001000001100101100111100",
						 "001000001100101010100110",
						 "001000001100101000010000",
						 "001000001100100101111010",
						 "001000001100100011100100",
						 "001000001101000110111101",
						 "001000001101000100100110",
						 "001000001101000010001111",
						 "001000001100111111111000",
						 "001000001100111101100001",
						 "001000001100111011001010",
						 "001000001100111000110011",
						 "001000001100110110011100",
						 "001000001100110100000101",
						 "001000001100110001101110",
						 "001000001100101111010111",
						 "001000001100101101000000",
						 "001000001100101010101001",
						 "001000001100101000010010",
						 "001000001100100101111011",
						 "001000001100100011100100",
						 "001000001010100011111111",
						 "001000001010100001101000",
						 "001000001010011111010001",
						 "001000001010011100111010",
						 "001000001010011010100011",
						 "001000001010011000001100",
						 "001000001010010101110101",
						 "001000001010010011011110",
						 "001000001010010001000111",
						 "001000001010001110110000",
						 "001000001010001100011001",
						 "001000001010001010000010",
						 "001000001010000111101011",
						 "001000001010000101010100",
						 "001000001010000010111101",
						 "001000001010000000100110",
						 "001000001010100011111111",
						 "001000001010100001101000",
						 "001000001010011111010001",
						 "001000001010011100111010",
						 "001000001010011010100011",
						 "001000001010011000001100",
						 "001000001010010101110101",
						 "001000001010010011011110",
						 "001000001010010001000111",
						 "001000001010001110110000",
						 "001000001010001100011001",
						 "001000001010001010000010",
						 "001000001010000111101011",
						 "001000001010000101010100",
						 "001000001010000010111101",
						 "001000001010000000100110",
						 "001000001010100100001110",
						 "001000001010100001110110",
						 "001000001010011111011110",
						 "001000001010011101000110",
						 "001000001010011010101110",
						 "001000001010011000010110",
						 "001000001010010101111110",
						 "001000001010010011100110",
						 "001000001010010001001110",
						 "001000001010001110110110",
						 "001000001010001100011110",
						 "001000001010001010000110",
						 "001000001010000111101110",
						 "001000001010000101010110",
						 "001000001010000010111110",
						 "001000001010000000100110",
						 "001000001010100100001110",
						 "001000001010100001110110",
						 "001000001010011111011110",
						 "001000001010011101000110",
						 "001000001010011010101110",
						 "001000001010011000010110",
						 "001000001010010101111110",
						 "001000001010010011100110",
						 "001000001010010001001110",
						 "001000001010001110110110",
						 "001000001010001100011110",
						 "001000001010001010000110",
						 "001000001010000111101110",
						 "001000001010000101010110",
						 "001000001010000010111110",
						 "001000001010000000100110",
						 "001000001000000001010000",
						 "001000000111111110111000",
						 "001000000111111100100000",
						 "001000000111111010001000",
						 "001000000111110111110000",
						 "001000000111110101011000",
						 "001000000111110011000000",
						 "001000000111110000101000",
						 "001000000111101110010000",
						 "001000000111101011111000",
						 "001000000111101001100000",
						 "001000000111100111001000",
						 "001000000111100100110000",
						 "001000000111100010011000",
						 "001000000111100000000000",
						 "001000000111011101101000",
						 "001000001000000001011111",
						 "001000000111111111000110",
						 "001000000111111100101101",
						 "001000000111111010010100",
						 "001000000111110111111011",
						 "001000000111110101100010",
						 "001000000111110011001001",
						 "001000000111110000110000",
						 "001000000111101110010111",
						 "001000000111101011111110",
						 "001000000111101001100101",
						 "001000000111100111001100",
						 "001000000111100100110011",
						 "001000000111100010011010",
						 "001000000111100000000001",
						 "001000000111011101101000",
						 "001000001000000001011111",
						 "001000000111111111000110",
						 "001000000111111100101101",
						 "001000000111111010010100",
						 "001000000111110111111011",
						 "001000000111110101100010",
						 "001000000111110011001001",
						 "001000000111110000110000",
						 "001000000111101110010111",
						 "001000000111101011111110",
						 "001000000111101001100101",
						 "001000000111100111001100",
						 "001000000111100100110011",
						 "001000000111100010011010",
						 "001000000111100000000001",
						 "001000000111011101101000",
						 "001000001000000001011111",
						 "001000000111111111000110",
						 "001000000111111100101101",
						 "001000000111111010010100",
						 "001000000111110111111011",
						 "001000000111110101100010",
						 "001000000111110011001001",
						 "001000000111110000110000",
						 "001000000111101110010111",
						 "001000000111101011111110",
						 "001000000111101001100101",
						 "001000000111100111001100",
						 "001000000111100100110011",
						 "001000000111100010011010",
						 "001000000111100000000001",
						 "001000000111011101101000",
						 "001000000101011110110000",
						 "001000000101011100010110",
						 "001000000101011001111100",
						 "001000000101010111100010",
						 "001000000101010101001000",
						 "001000000101010010101110",
						 "001000000101010000010100",
						 "001000000101001101111010",
						 "001000000101001011100000",
						 "001000000101001001000110",
						 "001000000101000110101100",
						 "001000000101000100010010",
						 "001000000101000001111000",
						 "001000000100111111011110",
						 "001000000100111101000100",
						 "001000000100111010101010",
						 "001000000101011110110000",
						 "001000000101011100010110",
						 "001000000101011001111100",
						 "001000000101010111100010",
						 "001000000101010101001000",
						 "001000000101010010101110",
						 "001000000101010000010100",
						 "001000000101001101111010",
						 "001000000101001011100000",
						 "001000000101001001000110",
						 "001000000101000110101100",
						 "001000000101000100010010",
						 "001000000101000001111000",
						 "001000000100111111011110",
						 "001000000100111101000100",
						 "001000000100111010101010",
						 "001000000101011110110000",
						 "001000000101011100010110",
						 "001000000101011001111100",
						 "001000000101010111100010",
						 "001000000101010101001000",
						 "001000000101010010101110",
						 "001000000101010000010100",
						 "001000000101001101111010",
						 "001000000101001011100000",
						 "001000000101001001000110",
						 "001000000101000110101100",
						 "001000000101000100010010",
						 "001000000101000001111000",
						 "001000000100111111011110",
						 "001000000100111101000100",
						 "001000000100111010101010",
						 "001000000101011110111111",
						 "001000000101011100100100",
						 "001000000101011010001001",
						 "001000000101010111101110",
						 "001000000101010101010011",
						 "001000000101010010111000",
						 "001000000101010000011101",
						 "001000000101001110000010",
						 "001000000101001011100111",
						 "001000000101001001001100",
						 "001000000101000110110001",
						 "001000000101000100010110",
						 "001000000101000001111011",
						 "001000000100111111100000",
						 "001000000100111101000101",
						 "001000000100111010101010",
						 "001000000010111100000001",
						 "001000000010111001100110",
						 "001000000010110111001011",
						 "001000000010110100110000",
						 "001000000010110010010101",
						 "001000000010101111111010",
						 "001000000010101101011111",
						 "001000000010101011000100",
						 "001000000010101000101001",
						 "001000000010100110001110",
						 "001000000010100011110011",
						 "001000000010100001011000",
						 "001000000010011110111101",
						 "001000000010011100100010",
						 "001000000010011010000111",
						 "001000000010010111101100",
						 "001000000010111100000001",
						 "001000000010111001100110",
						 "001000000010110111001011",
						 "001000000010110100110000",
						 "001000000010110010010101",
						 "001000000010101111111010",
						 "001000000010101101011111",
						 "001000000010101011000100",
						 "001000000010101000101001",
						 "001000000010100110001110",
						 "001000000010100011110011",
						 "001000000010100001011000",
						 "001000000010011110111101",
						 "001000000010011100100010",
						 "001000000010011010000111",
						 "001000000010010111101100",
						 "001000000010111100000001",
						 "001000000010111001100110",
						 "001000000010110111001011",
						 "001000000010110100110000",
						 "001000000010110010010101",
						 "001000000010101111111010",
						 "001000000010101101011111",
						 "001000000010101011000100",
						 "001000000010101000101001",
						 "001000000010100110001110",
						 "001000000010100011110011",
						 "001000000010100001011000",
						 "001000000010011110111101",
						 "001000000010011100100010",
						 "001000000010011010000111",
						 "001000000010010111101100",
						 "001000000010111100010000",
						 "001000000010111001110100",
						 "001000000010110111011000",
						 "001000000010110100111100",
						 "001000000010110010100000",
						 "001000000010110000000100",
						 "001000000010101101101000",
						 "001000000010101011001100",
						 "001000000010101000110000",
						 "001000000010100110010100",
						 "001000000010100011111000",
						 "001000000010100001011100",
						 "001000000010011111000000",
						 "001000000010011100100100",
						 "001000000010011010001000",
						 "001000000010010111101100",
						 "001000000010111100010000",
						 "001000000010111001110100",
						 "001000000010110111011000",
						 "001000000010110100111100",
						 "001000000010110010100000",
						 "001000000010110000000100",
						 "001000000010101101101000",
						 "001000000010101011001100",
						 "001000000010101000110000",
						 "001000000010100110010100",
						 "001000000010100011111000",
						 "001000000010100001011100",
						 "001000000010011111000000",
						 "001000000010011100100100",
						 "001000000010011010001000",
						 "001000000010010111101100",
						 "001000000000011001010010",
						 "001000000000010110110110",
						 "001000000000010100011010",
						 "001000000000010001111110",
						 "001000000000001111100010",
						 "001000000000001101000110",
						 "001000000000001010101010",
						 "001000000000001000001110",
						 "001000000000000101110010",
						 "001000000000000011010110",
						 "001000000000000000111010",
						 "000111111111111110011110",
						 "000111111111111100000010",
						 "000111111111111001100110",
						 "000111111111110111001010",
						 "000111111111110100101110",
						 "001000000000011001100001",
						 "001000000000010111000100",
						 "001000000000010100100111",
						 "001000000000010010001010",
						 "001000000000001111101101",
						 "001000000000001101010000",
						 "001000000000001010110011",
						 "001000000000001000010110",
						 "001000000000000101111001",
						 "001000000000000011011100",
						 "001000000000000000111111",
						 "000111111111111110100010",
						 "000111111111111100000101",
						 "000111111111111001101000",
						 "000111111111110111001011",
						 "000111111111110100101110",
						 "001000000000011001100001",
						 "001000000000010111000100",
						 "001000000000010100100111",
						 "001000000000010010001010",
						 "001000000000001111101101",
						 "001000000000001101010000",
						 "001000000000001010110011",
						 "001000000000001000010110",
						 "001000000000000101111001",
						 "001000000000000011011100",
						 "001000000000000000111111",
						 "000111111111111110100010",
						 "000111111111111100000101",
						 "000111111111111001101000",
						 "000111111111110111001011",
						 "000111111111110100101110",
						 "001000000000011001100001",
						 "001000000000010111000100",
						 "001000000000010100100111",
						 "001000000000010010001010",
						 "001000000000001111101101",
						 "001000000000001101010000",
						 "001000000000001010110011",
						 "001000000000001000010110",
						 "001000000000000101111001",
						 "001000000000000011011100",
						 "001000000000000000111111",
						 "000111111111111110100010",
						 "000111111111111100000101",
						 "000111111111111001101000",
						 "000111111111110111001011",
						 "000111111111110100101110",
						 "000111111101110110110010",
						 "000111111101110100010100",
						 "000111111101110001110110",
						 "000111111101101111011000",
						 "000111111101101100111010",
						 "000111111101101010011100",
						 "000111111101100111111110",
						 "000111111101100101100000",
						 "000111111101100011000010",
						 "000111111101100000100100",
						 "000111111101011110000110",
						 "000111111101011011101000",
						 "000111111101011001001010",
						 "000111111101010110101100",
						 "000111111101010100001110",
						 "000111111101010001110000",
						 "000111111101110110110010",
						 "000111111101110100010100",
						 "000111111101110001110110",
						 "000111111101101111011000",
						 "000111111101101100111010",
						 "000111111101101010011100",
						 "000111111101100111111110",
						 "000111111101100101100000",
						 "000111111101100011000010",
						 "000111111101100000100100",
						 "000111111101011110000110",
						 "000111111101011011101000",
						 "000111111101011001001010",
						 "000111111101010110101100",
						 "000111111101010100001110",
						 "000111111101010001110000",
						 "000111111101110110110010",
						 "000111111101110100010100",
						 "000111111101110001110110",
						 "000111111101101111011000",
						 "000111111101101100111010",
						 "000111111101101010011100",
						 "000111111101100111111110",
						 "000111111101100101100000",
						 "000111111101100011000010",
						 "000111111101100000100100",
						 "000111111101011110000110",
						 "000111111101011011101000",
						 "000111111101011001001010",
						 "000111111101010110101100",
						 "000111111101010100001110",
						 "000111111101010001110000",
						 "000111111101110111000001",
						 "000111111101110100100010",
						 "000111111101110010000011",
						 "000111111101101111100100",
						 "000111111101101101000101",
						 "000111111101101010100110",
						 "000111111101101000000111",
						 "000111111101100101101000",
						 "000111111101100011001001",
						 "000111111101100000101010",
						 "000111111101011110001011",
						 "000111111101011011101100",
						 "000111111101011001001101",
						 "000111111101010110101110",
						 "000111111101010100001111",
						 "000111111101010001110000",
						 "000111111011010100000011",
						 "000111111011010001100100",
						 "000111111011001111000101",
						 "000111111011001100100110",
						 "000111111011001010000111",
						 "000111111011000111101000",
						 "000111111011000101001001",
						 "000111111011000010101010",
						 "000111111011000000001011",
						 "000111111010111101101100",
						 "000111111010111011001101",
						 "000111111010111000101110",
						 "000111111010110110001111",
						 "000111111010110011110000",
						 "000111111010110001010001",
						 "000111111010101110110010",
						 "000111111011010100000011",
						 "000111111011010001100100",
						 "000111111011001111000101",
						 "000111111011001100100110",
						 "000111111011001010000111",
						 "000111111011000111101000",
						 "000111111011000101001001",
						 "000111111011000010101010",
						 "000111111011000000001011",
						 "000111111010111101101100",
						 "000111111010111011001101",
						 "000111111010111000101110",
						 "000111111010110110001111",
						 "000111111010110011110000",
						 "000111111010110001010001",
						 "000111111010101110110010",
						 "000111111011010100000011",
						 "000111111011010001100100",
						 "000111111011001111000101",
						 "000111111011001100100110",
						 "000111111011001010000111",
						 "000111111011000111101000",
						 "000111111011000101001001",
						 "000111111011000010101010",
						 "000111111011000000001011",
						 "000111111010111101101100",
						 "000111111010111011001101",
						 "000111111010111000101110",
						 "000111111010110110001111",
						 "000111111010110011110000",
						 "000111111010110001010001",
						 "000111111010101110110010",
						 "000111111011010100010010",
						 "000111111011010001110010",
						 "000111111011001111010010",
						 "000111111011001100110010",
						 "000111111011001010010010",
						 "000111111011000111110010",
						 "000111111011000101010010",
						 "000111111011000010110010",
						 "000111111011000000010010",
						 "000111111010111101110010",
						 "000111111010111011010010",
						 "000111111010111000110010",
						 "000111111010110110010010",
						 "000111111010110011110010",
						 "000111111010110001010010",
						 "000111111010101110110010",
						 "000111111000110001010100",
						 "000111111000101110110100",
						 "000111111000101100010100",
						 "000111111000101001110100",
						 "000111111000100111010100",
						 "000111111000100100110100",
						 "000111111000100010010100",
						 "000111111000011111110100",
						 "000111111000011101010100",
						 "000111111000011010110100",
						 "000111111000011000010100",
						 "000111111000010101110100",
						 "000111111000010011010100",
						 "000111111000010000110100",
						 "000111111000001110010100",
						 "000111111000001011110100",
						 "000111111000110001010100",
						 "000111111000101110110100",
						 "000111111000101100010100",
						 "000111111000101001110100",
						 "000111111000100111010100",
						 "000111111000100100110100",
						 "000111111000100010010100",
						 "000111111000011111110100",
						 "000111111000011101010100",
						 "000111111000011010110100",
						 "000111111000011000010100",
						 "000111111000010101110100",
						 "000111111000010011010100",
						 "000111111000010000110100",
						 "000111111000001110010100",
						 "000111111000001011110100",
						 "000111111000110001100011",
						 "000111111000101111000010",
						 "000111111000101100100001",
						 "000111111000101010000000",
						 "000111111000100111011111",
						 "000111111000100100111110",
						 "000111111000100010011101",
						 "000111111000011111111100",
						 "000111111000011101011011",
						 "000111111000011010111010",
						 "000111111000011000011001",
						 "000111111000010101111000",
						 "000111111000010011010111",
						 "000111111000010000110110",
						 "000111111000001110010101",
						 "000111111000001011110100",
						 "000111111000110001100011",
						 "000111111000101111000010",
						 "000111111000101100100001",
						 "000111111000101010000000",
						 "000111111000100111011111",
						 "000111111000100100111110",
						 "000111111000100010011101",
						 "000111111000011111111100",
						 "000111111000011101011011",
						 "000111111000011010111010",
						 "000111111000011000011001",
						 "000111111000010101111000",
						 "000111111000010011010111",
						 "000111111000010000110110",
						 "000111111000001110010101",
						 "000111111000001011110100",
						 "000111110110001110100101",
						 "000111110110001100000100",
						 "000111110110001001100011",
						 "000111110110000111000010",
						 "000111110110000100100001",
						 "000111110110000010000000",
						 "000111110101111111011111",
						 "000111110101111100111110",
						 "000111110101111010011101",
						 "000111110101110111111100",
						 "000111110101110101011011",
						 "000111110101110010111010",
						 "000111110101110000011001",
						 "000111110101101101111000",
						 "000111110101101011010111",
						 "000111110101101000110110",
						 "000111110110001110110100",
						 "000111110110001100010010",
						 "000111110110001001110000",
						 "000111110110000111001110",
						 "000111110110000100101100",
						 "000111110110000010001010",
						 "000111110101111111101000",
						 "000111110101111101000110",
						 "000111110101111010100100",
						 "000111110101111000000010",
						 "000111110101110101100000",
						 "000111110101110010111110",
						 "000111110101110000011100",
						 "000111110101101101111010",
						 "000111110101101011011000",
						 "000111110101101000110110",
						 "000111110110001110110100",
						 "000111110110001100010010",
						 "000111110110001001110000",
						 "000111110110000111001110",
						 "000111110110000100101100",
						 "000111110110000010001010",
						 "000111110101111111101000",
						 "000111110101111101000110",
						 "000111110101111010100100",
						 "000111110101111000000010",
						 "000111110101110101100000",
						 "000111110101110010111110",
						 "000111110101110000011100",
						 "000111110101101101111010",
						 "000111110101101011011000",
						 "000111110101101000110110",
						 "000111110110001110110100",
						 "000111110110001100010010",
						 "000111110110001001110000",
						 "000111110110000111001110",
						 "000111110110000100101100",
						 "000111110110000010001010",
						 "000111110101111111101000",
						 "000111110101111101000110",
						 "000111110101111010100100",
						 "000111110101111000000010",
						 "000111110101110101100000",
						 "000111110101110010111110",
						 "000111110101110000011100",
						 "000111110101101101111010",
						 "000111110101101011011000",
						 "000111110101101000110110",
						 "000111110011101100000101",
						 "000111110011101001100010",
						 "000111110011100110111111",
						 "000111110011100100011100",
						 "000111110011100001111001",
						 "000111110011011111010110",
						 "000111110011011100110011",
						 "000111110011011010010000",
						 "000111110011010111101101",
						 "000111110011010101001010",
						 "000111110011010010100111",
						 "000111110011010000000100",
						 "000111110011001101100001",
						 "000111110011001010111110",
						 "000111110011001000011011",
						 "000111110011000101111000",
						 "000111110011101100000101",
						 "000111110011101001100010",
						 "000111110011100110111111",
						 "000111110011100100011100",
						 "000111110011100001111001",
						 "000111110011011111010110",
						 "000111110011011100110011",
						 "000111110011011010010000",
						 "000111110011010111101101",
						 "000111110011010101001010",
						 "000111110011010010100111",
						 "000111110011010000000100",
						 "000111110011001101100001",
						 "000111110011001010111110",
						 "000111110011001000011011",
						 "000111110011000101111000",
						 "000111110011101100000101",
						 "000111110011101001100010",
						 "000111110011100110111111",
						 "000111110011100100011100",
						 "000111110011100001111001",
						 "000111110011011111010110",
						 "000111110011011100110011",
						 "000111110011011010010000",
						 "000111110011010111101101",
						 "000111110011010101001010",
						 "000111110011010010100111",
						 "000111110011010000000100",
						 "000111110011001101100001",
						 "000111110011001010111110",
						 "000111110011001000011011",
						 "000111110011000101111000",
						 "000111110011101100000101",
						 "000111110011101001100010",
						 "000111110011100110111111",
						 "000111110011100100011100",
						 "000111110011100001111001",
						 "000111110011011111010110",
						 "000111110011011100110011",
						 "000111110011011010010000",
						 "000111110011010111101101",
						 "000111110011010101001010",
						 "000111110011010010100111",
						 "000111110011010000000100",
						 "000111110011001101100001",
						 "000111110011001010111110",
						 "000111110011001000011011",
						 "000111110011000101111000",
						 "000111110001001001010110",
						 "000111110001000110110010",
						 "000111110001000100001110",
						 "000111110001000001101010",
						 "000111110000111111000110",
						 "000111110000111100100010",
						 "000111110000111001111110",
						 "000111110000110111011010",
						 "000111110000110100110110",
						 "000111110000110010010010",
						 "000111110000101111101110",
						 "000111110000101101001010",
						 "000111110000101010100110",
						 "000111110000101000000010",
						 "000111110000100101011110",
						 "000111110000100010111010",
						 "000111110001001001010110",
						 "000111110001000110110010",
						 "000111110001000100001110",
						 "000111110001000001101010",
						 "000111110000111111000110",
						 "000111110000111100100010",
						 "000111110000111001111110",
						 "000111110000110111011010",
						 "000111110000110100110110",
						 "000111110000110010010010",
						 "000111110000101111101110",
						 "000111110000101101001010",
						 "000111110000101010100110",
						 "000111110000101000000010",
						 "000111110000100101011110",
						 "000111110000100010111010",
						 "000111110001001001010110",
						 "000111110001000110110010",
						 "000111110001000100001110",
						 "000111110001000001101010",
						 "000111110000111111000110",
						 "000111110000111100100010",
						 "000111110000111001111110",
						 "000111110000110111011010",
						 "000111110000110100110110",
						 "000111110000110010010010",
						 "000111110000101111101110",
						 "000111110000101101001010",
						 "000111110000101010100110",
						 "000111110000101000000010",
						 "000111110000100101011110",
						 "000111110000100010111010",
						 "000111110001001001100101",
						 "000111110001000111000000",
						 "000111110001000100011011",
						 "000111110001000001110110",
						 "000111110000111111010001",
						 "000111110000111100101100",
						 "000111110000111010000111",
						 "000111110000110111100010",
						 "000111110000110100111101",
						 "000111110000110010011000",
						 "000111110000101111110011",
						 "000111110000101101001110",
						 "000111110000101010101001",
						 "000111110000101000000100",
						 "000111110000100101011111",
						 "000111110000100010111010",
						 "000111101110100110100111",
						 "000111101110100100000010",
						 "000111101110100001011101",
						 "000111101110011110111000",
						 "000111101110011100010011",
						 "000111101110011001101110",
						 "000111101110010111001001",
						 "000111101110010100100100",
						 "000111101110010001111111",
						 "000111101110001111011010",
						 "000111101110001100110101",
						 "000111101110001010010000",
						 "000111101110000111101011",
						 "000111101110000101000110",
						 "000111101110000010100001",
						 "000111101101111111111100",
						 "000111101110100110100111",
						 "000111101110100100000010",
						 "000111101110100001011101",
						 "000111101110011110111000",
						 "000111101110011100010011",
						 "000111101110011001101110",
						 "000111101110010111001001",
						 "000111101110010100100100",
						 "000111101110010001111111",
						 "000111101110001111011010",
						 "000111101110001100110101",
						 "000111101110001010010000",
						 "000111101110000111101011",
						 "000111101110000101000110",
						 "000111101110000010100001",
						 "000111101101111111111100",
						 "000111101110100110110110",
						 "000111101110100100010000",
						 "000111101110100001101010",
						 "000111101110011111000100",
						 "000111101110011100011110",
						 "000111101110011001111000",
						 "000111101110010111010010",
						 "000111101110010100101100",
						 "000111101110010010000110",
						 "000111101110001111100000",
						 "000111101110001100111010",
						 "000111101110001010010100",
						 "000111101110000111101110",
						 "000111101110000101001000",
						 "000111101110000010100010",
						 "000111101101111111111100",
						 "000111101110100110110110",
						 "000111101110100100010000",
						 "000111101110100001101010",
						 "000111101110011111000100",
						 "000111101110011100011110",
						 "000111101110011001111000",
						 "000111101110010111010010",
						 "000111101110010100101100",
						 "000111101110010010000110",
						 "000111101110001111100000",
						 "000111101110001100111010",
						 "000111101110001010010100",
						 "000111101110000111101110",
						 "000111101110000101001000",
						 "000111101110000010100010",
						 "000111101101111111111100",
						 "000111101100000011111000",
						 "000111101100000001010010",
						 "000111101011111110101100",
						 "000111101011111100000110",
						 "000111101011111001100000",
						 "000111101011110110111010",
						 "000111101011110100010100",
						 "000111101011110001101110",
						 "000111101011101111001000",
						 "000111101011101100100010",
						 "000111101011101001111100",
						 "000111101011100111010110",
						 "000111101011100100110000",
						 "000111101011100010001010",
						 "000111101011011111100100",
						 "000111101011011100111110",
						 "000111101100000011111000",
						 "000111101100000001010010",
						 "000111101011111110101100",
						 "000111101011111100000110",
						 "000111101011111001100000",
						 "000111101011110110111010",
						 "000111101011110100010100",
						 "000111101011110001101110",
						 "000111101011101111001000",
						 "000111101011101100100010",
						 "000111101011101001111100",
						 "000111101011100111010110",
						 "000111101011100100110000",
						 "000111101011100010001010",
						 "000111101011011111100100",
						 "000111101011011100111110",
						 "000111101100000100000111",
						 "000111101100000001100000",
						 "000111101011111110111001",
						 "000111101011111100010010",
						 "000111101011111001101011",
						 "000111101011110111000100",
						 "000111101011110100011101",
						 "000111101011110001110110",
						 "000111101011101111001111",
						 "000111101011101100101000",
						 "000111101011101010000001",
						 "000111101011100111011010",
						 "000111101011100100110011",
						 "000111101011100010001100",
						 "000111101011011111100101",
						 "000111101011011100111110",
						 "000111101100000100000111",
						 "000111101100000001100000",
						 "000111101011111110111001",
						 "000111101011111100010010",
						 "000111101011111001101011",
						 "000111101011110111000100",
						 "000111101011110100011101",
						 "000111101011110001110110",
						 "000111101011101111001111",
						 "000111101011101100101000",
						 "000111101011101010000001",
						 "000111101011100111011010",
						 "000111101011100100110011",
						 "000111101011100010001100",
						 "000111101011011111100101",
						 "000111101011011100111110",
						 "000111101001100001001001",
						 "000111101001011110100010",
						 "000111101001011011111011",
						 "000111101001011001010100",
						 "000111101001010110101101",
						 "000111101001010100000110",
						 "000111101001010001011111",
						 "000111101001001110111000",
						 "000111101001001100010001",
						 "000111101001001001101010",
						 "000111101001000111000011",
						 "000111101001000100011100",
						 "000111101001000001110101",
						 "000111101000111111001110",
						 "000111101000111100100111",
						 "000111101000111010000000",
						 "000111101001100001011000",
						 "000111101001011110110000",
						 "000111101001011100001000",
						 "000111101001011001100000",
						 "000111101001010110111000",
						 "000111101001010100010000",
						 "000111101001010001101000",
						 "000111101001001111000000",
						 "000111101001001100011000",
						 "000111101001001001110000",
						 "000111101001000111001000",
						 "000111101001000100100000",
						 "000111101001000001111000",
						 "000111101000111111010000",
						 "000111101000111100101000",
						 "000111101000111010000000",
						 "000111101001100001011000",
						 "000111101001011110110000",
						 "000111101001011100001000",
						 "000111101001011001100000",
						 "000111101001010110111000",
						 "000111101001010100010000",
						 "000111101001010001101000",
						 "000111101001001111000000",
						 "000111101001001100011000",
						 "000111101001001001110000",
						 "000111101001000111001000",
						 "000111101001000100100000",
						 "000111101001000001111000",
						 "000111101000111111010000",
						 "000111101000111100101000",
						 "000111101000111010000000",
						 "000111101001100001011000",
						 "000111101001011110110000",
						 "000111101001011100001000",
						 "000111101001011001100000",
						 "000111101001010110111000",
						 "000111101001010100010000",
						 "000111101001010001101000",
						 "000111101001001111000000",
						 "000111101001001100011000",
						 "000111101001001001110000",
						 "000111101001000111001000",
						 "000111101001000100100000",
						 "000111101001000001111000",
						 "000111101000111111010000",
						 "000111101000111100101000",
						 "000111101000111010000000",
						 "000111100110111110011010",
						 "000111100110111011110010",
						 "000111100110111001001010",
						 "000111100110110110100010",
						 "000111100110110011111010",
						 "000111100110110001010010",
						 "000111100110101110101010",
						 "000111100110101100000010",
						 "000111100110101001011010",
						 "000111100110100110110010",
						 "000111100110100100001010",
						 "000111100110100001100010",
						 "000111100110011110111010",
						 "000111100110011100010010",
						 "000111100110011001101010",
						 "000111100110010111000010",
						 "000111100110111110101001",
						 "000111100110111100000000",
						 "000111100110111001010111",
						 "000111100110110110101110",
						 "000111100110110100000101",
						 "000111100110110001011100",
						 "000111100110101110110011",
						 "000111100110101100001010",
						 "000111100110101001100001",
						 "000111100110100110111000",
						 "000111100110100100001111",
						 "000111100110100001100110",
						 "000111100110011110111101",
						 "000111100110011100010100",
						 "000111100110011001101011",
						 "000111100110010111000010",
						 "000111100110111110101001",
						 "000111100110111100000000",
						 "000111100110111001010111",
						 "000111100110110110101110",
						 "000111100110110100000101",
						 "000111100110110001011100",
						 "000111100110101110110011",
						 "000111100110101100001010",
						 "000111100110101001100001",
						 "000111100110100110111000",
						 "000111100110100100001111",
						 "000111100110100001100110",
						 "000111100110011110111101",
						 "000111100110011100010100",
						 "000111100110011001101011",
						 "000111100110010111000010",
						 "000111100110111110101001",
						 "000111100110111100000000",
						 "000111100110111001010111",
						 "000111100110110110101110",
						 "000111100110110100000101",
						 "000111100110110001011100",
						 "000111100110101110110011",
						 "000111100110101100001010",
						 "000111100110101001100001",
						 "000111100110100110111000",
						 "000111100110100100001111",
						 "000111100110100001100110",
						 "000111100110011110111101",
						 "000111100110011100010100",
						 "000111100110011001101011",
						 "000111100110010111000010",
						 "000111100100011011111010",
						 "000111100100011001010000",
						 "000111100100010110100110",
						 "000111100100010011111100",
						 "000111100100010001010010",
						 "000111100100001110101000",
						 "000111100100001011111110",
						 "000111100100001001010100",
						 "000111100100000110101010",
						 "000111100100000100000000",
						 "000111100100000001010110",
						 "000111100011111110101100",
						 "000111100011111100000010",
						 "000111100011111001011000",
						 "000111100011110110101110",
						 "000111100011110100000100",
						 "000111100100011011111010",
						 "000111100100011001010000",
						 "000111100100010110100110",
						 "000111100100010011111100",
						 "000111100100010001010010",
						 "000111100100001110101000",
						 "000111100100001011111110",
						 "000111100100001001010100",
						 "000111100100000110101010",
						 "000111100100000100000000",
						 "000111100100000001010110",
						 "000111100011111110101100",
						 "000111100011111100000010",
						 "000111100011111001011000",
						 "000111100011110110101110",
						 "000111100011110100000100",
						 "000111100100011011111010",
						 "000111100100011001010000",
						 "000111100100010110100110",
						 "000111100100010011111100",
						 "000111100100010001010010",
						 "000111100100001110101000",
						 "000111100100001011111110",
						 "000111100100001001010100",
						 "000111100100000110101010",
						 "000111100100000100000000",
						 "000111100100000001010110",
						 "000111100011111110101100",
						 "000111100011111100000010",
						 "000111100011111001011000",
						 "000111100011110110101110",
						 "000111100011110100000100",
						 "000111100001111001001011",
						 "000111100001110110100000",
						 "000111100001110011110101",
						 "000111100001110001001010",
						 "000111100001101110011111",
						 "000111100001101011110100",
						 "000111100001101001001001",
						 "000111100001100110011110",
						 "000111100001100011110011",
						 "000111100001100001001000",
						 "000111100001011110011101",
						 "000111100001011011110010",
						 "000111100001011001000111",
						 "000111100001010110011100",
						 "000111100001010011110001",
						 "000111100001010001000110",
						 "000111100001111001001011",
						 "000111100001110110100000",
						 "000111100001110011110101",
						 "000111100001110001001010",
						 "000111100001101110011111",
						 "000111100001101011110100",
						 "000111100001101001001001",
						 "000111100001100110011110",
						 "000111100001100011110011",
						 "000111100001100001001000",
						 "000111100001011110011101",
						 "000111100001011011110010",
						 "000111100001011001000111",
						 "000111100001010110011100",
						 "000111100001010011110001",
						 "000111100001010001000110",
						 "000111100001111001001011",
						 "000111100001110110100000",
						 "000111100001110011110101",
						 "000111100001110001001010",
						 "000111100001101110011111",
						 "000111100001101011110100",
						 "000111100001101001001001",
						 "000111100001100110011110",
						 "000111100001100011110011",
						 "000111100001100001001000",
						 "000111100001011110011101",
						 "000111100001011011110010",
						 "000111100001011001000111",
						 "000111100001010110011100",
						 "000111100001010011110001",
						 "000111100001010001000110",
						 "000111100001111001001011",
						 "000111100001110110100000",
						 "000111100001110011110101",
						 "000111100001110001001010",
						 "000111100001101110011111",
						 "000111100001101011110100",
						 "000111100001101001001001",
						 "000111100001100110011110",
						 "000111100001100011110011",
						 "000111100001100001001000",
						 "000111100001011110011101",
						 "000111100001011011110010",
						 "000111100001011001000111",
						 "000111100001010110011100",
						 "000111100001010011110001",
						 "000111100001010001000110",
						 "000111011111010110011100",
						 "000111011111010011110000",
						 "000111011111010001000100",
						 "000111011111001110011000",
						 "000111011111001011101100",
						 "000111011111001001000000",
						 "000111011111000110010100",
						 "000111011111000011101000",
						 "000111011111000000111100",
						 "000111011110111110010000",
						 "000111011110111011100100",
						 "000111011110111000111000",
						 "000111011110110110001100",
						 "000111011110110011100000",
						 "000111011110110000110100",
						 "000111011110101110001000",
						 "000111011111010110011100",
						 "000111011111010011110000",
						 "000111011111010001000100",
						 "000111011111001110011000",
						 "000111011111001011101100",
						 "000111011111001001000000",
						 "000111011111000110010100",
						 "000111011111000011101000",
						 "000111011111000000111100",
						 "000111011110111110010000",
						 "000111011110111011100100",
						 "000111011110111000111000",
						 "000111011110110110001100",
						 "000111011110110011100000",
						 "000111011110110000110100",
						 "000111011110101110001000",
						 "000111011111010110011100",
						 "000111011111010011110000",
						 "000111011111010001000100",
						 "000111011111001110011000",
						 "000111011111001011101100",
						 "000111011111001001000000",
						 "000111011111000110010100",
						 "000111011111000011101000",
						 "000111011111000000111100",
						 "000111011110111110010000",
						 "000111011110111011100100",
						 "000111011110111000111000",
						 "000111011110110110001100",
						 "000111011110110011100000",
						 "000111011110110000110100",
						 "000111011110101110001000",
						 "000111011111010110101011",
						 "000111011111010011111110",
						 "000111011111010001010001",
						 "000111011111001110100100",
						 "000111011111001011110111",
						 "000111011111001001001010",
						 "000111011111000110011101",
						 "000111011111000011110000",
						 "000111011111000001000011",
						 "000111011110111110010110",
						 "000111011110111011101001",
						 "000111011110111000111100",
						 "000111011110110110001111",
						 "000111011110110011100010",
						 "000111011110110000110101",
						 "000111011110101110001000",
						 "000111011100110011101101",
						 "000111011100110001000000",
						 "000111011100101110010011",
						 "000111011100101011100110",
						 "000111011100101000111001",
						 "000111011100100110001100",
						 "000111011100100011011111",
						 "000111011100100000110010",
						 "000111011100011110000101",
						 "000111011100011011011000",
						 "000111011100011000101011",
						 "000111011100010101111110",
						 "000111011100010011010001",
						 "000111011100010000100100",
						 "000111011100001101110111",
						 "000111011100001011001010",
						 "000111011100110011101101",
						 "000111011100110001000000",
						 "000111011100101110010011",
						 "000111011100101011100110",
						 "000111011100101000111001",
						 "000111011100100110001100",
						 "000111011100100011011111",
						 "000111011100100000110010",
						 "000111011100011110000101",
						 "000111011100011011011000",
						 "000111011100011000101011",
						 "000111011100010101111110",
						 "000111011100010011010001",
						 "000111011100010000100100",
						 "000111011100001101110111",
						 "000111011100001011001010",
						 "000111011100110011101101",
						 "000111011100110001000000",
						 "000111011100101110010011",
						 "000111011100101011100110",
						 "000111011100101000111001",
						 "000111011100100110001100",
						 "000111011100100011011111",
						 "000111011100100000110010",
						 "000111011100011110000101",
						 "000111011100011011011000",
						 "000111011100011000101011",
						 "000111011100010101111110",
						 "000111011100010011010001",
						 "000111011100010000100100",
						 "000111011100001101110111",
						 "000111011100001011001010",
						 "000111011100110011111100",
						 "000111011100110001001110",
						 "000111011100101110100000",
						 "000111011100101011110010",
						 "000111011100101001000100",
						 "000111011100100110010110",
						 "000111011100100011101000",
						 "000111011100100000111010",
						 "000111011100011110001100",
						 "000111011100011011011110",
						 "000111011100011000110000",
						 "000111011100010110000010",
						 "000111011100010011010100",
						 "000111011100010000100110",
						 "000111011100001101111000",
						 "000111011100001011001010",
						 "000111011010010000111110",
						 "000111011010001110010000",
						 "000111011010001011100010",
						 "000111011010001000110100",
						 "000111011010000110000110",
						 "000111011010000011011000",
						 "000111011010000000101010",
						 "000111011001111101111100",
						 "000111011001111011001110",
						 "000111011001111000100000",
						 "000111011001110101110010",
						 "000111011001110011000100",
						 "000111011001110000010110",
						 "000111011001101101101000",
						 "000111011001101010111010",
						 "000111011001101000001100",
						 "000111011010010000111110",
						 "000111011010001110010000",
						 "000111011010001011100010",
						 "000111011010001000110100",
						 "000111011010000110000110",
						 "000111011010000011011000",
						 "000111011010000000101010",
						 "000111011001111101111100",
						 "000111011001111011001110",
						 "000111011001111000100000",
						 "000111011001110101110010",
						 "000111011001110011000100",
						 "000111011001110000010110",
						 "000111011001101101101000",
						 "000111011001101010111010",
						 "000111011001101000001100",
						 "000111011010010001001101",
						 "000111011010001110011110",
						 "000111011010001011101111",
						 "000111011010001001000000",
						 "000111011010000110010001",
						 "000111011010000011100010",
						 "000111011010000000110011",
						 "000111011001111110000100",
						 "000111011001111011010101",
						 "000111011001111000100110",
						 "000111011001110101110111",
						 "000111011001110011001000",
						 "000111011001110000011001",
						 "000111011001101101101010",
						 "000111011001101010111011",
						 "000111011001101000001100",
						 "000111010111101110001111",
						 "000111010111101011100000",
						 "000111010111101000110001",
						 "000111010111100110000010",
						 "000111010111100011010011",
						 "000111010111100000100100",
						 "000111010111011101110101",
						 "000111010111011011000110",
						 "000111010111011000010111",
						 "000111010111010101101000",
						 "000111010111010010111001",
						 "000111010111010000001010",
						 "000111010111001101011011",
						 "000111010111001010101100",
						 "000111010111000111111101",
						 "000111010111000101001110",
						 "000111010111101110001111",
						 "000111010111101011100000",
						 "000111010111101000110001",
						 "000111010111100110000010",
						 "000111010111100011010011",
						 "000111010111100000100100",
						 "000111010111011101110101",
						 "000111010111011011000110",
						 "000111010111011000010111",
						 "000111010111010101101000",
						 "000111010111010010111001",
						 "000111010111010000001010",
						 "000111010111001101011011",
						 "000111010111001010101100",
						 "000111010111000111111101",
						 "000111010111000101001110",
						 "000111010111101110001111",
						 "000111010111101011100000",
						 "000111010111101000110001",
						 "000111010111100110000010",
						 "000111010111100011010011",
						 "000111010111100000100100",
						 "000111010111011101110101",
						 "000111010111011011000110",
						 "000111010111011000010111",
						 "000111010111010101101000",
						 "000111010111010010111001",
						 "000111010111010000001010",
						 "000111010111001101011011",
						 "000111010111001010101100",
						 "000111010111000111111101",
						 "000111010111000101001110",
						 "000111010111101110011110",
						 "000111010111101011101110",
						 "000111010111101000111110",
						 "000111010111100110001110",
						 "000111010111100011011110",
						 "000111010111100000101110",
						 "000111010111011101111110",
						 "000111010111011011001110",
						 "000111010111011000011110",
						 "000111010111010101101110",
						 "000111010111010010111110",
						 "000111010111010000001110",
						 "000111010111001101011110",
						 "000111010111001010101110",
						 "000111010111000111111110",
						 "000111010111000101001110",
						 "000111010101001011100000",
						 "000111010101001000110000",
						 "000111010101000110000000",
						 "000111010101000011010000",
						 "000111010101000000100000",
						 "000111010100111101110000",
						 "000111010100111011000000",
						 "000111010100111000010000",
						 "000111010100110101100000",
						 "000111010100110010110000",
						 "000111010100110000000000",
						 "000111010100101101010000",
						 "000111010100101010100000",
						 "000111010100100111110000",
						 "000111010100100101000000",
						 "000111010100100010010000",
						 "000111010101001011100000",
						 "000111010101001000110000",
						 "000111010101000110000000",
						 "000111010101000011010000",
						 "000111010101000000100000",
						 "000111010100111101110000",
						 "000111010100111011000000",
						 "000111010100111000010000",
						 "000111010100110101100000",
						 "000111010100110010110000",
						 "000111010100110000000000",
						 "000111010100101101010000",
						 "000111010100101010100000",
						 "000111010100100111110000",
						 "000111010100100101000000",
						 "000111010100100010010000",
						 "000111010101001011101111",
						 "000111010101001000111110",
						 "000111010101000110001101",
						 "000111010101000011011100",
						 "000111010101000000101011",
						 "000111010100111101111010",
						 "000111010100111011001001",
						 "000111010100111000011000",
						 "000111010100110101100111",
						 "000111010100110010110110",
						 "000111010100110000000101",
						 "000111010100101101010100",
						 "000111010100101010100011",
						 "000111010100100111110010",
						 "000111010100100101000001",
						 "000111010100100010010000",
						 "000111010101001011101111",
						 "000111010101001000111110",
						 "000111010101000110001101",
						 "000111010101000011011100",
						 "000111010101000000101011",
						 "000111010100111101111010",
						 "000111010100111011001001",
						 "000111010100111000011000",
						 "000111010100110101100111",
						 "000111010100110010110110",
						 "000111010100110000000101",
						 "000111010100101101010100",
						 "000111010100101010100011",
						 "000111010100100111110010",
						 "000111010100100101000001",
						 "000111010100100010010000",
						 "000111010010101000110001",
						 "000111010010100110000000",
						 "000111010010100011001111",
						 "000111010010100000011110",
						 "000111010010011101101101",
						 "000111010010011010111100",
						 "000111010010011000001011",
						 "000111010010010101011010",
						 "000111010010010010101001",
						 "000111010010001111111000",
						 "000111010010001101000111",
						 "000111010010001010010110",
						 "000111010010000111100101",
						 "000111010010000100110100",
						 "000111010010000010000011",
						 "000111010001111111010010",
						 "000111010010101000110001",
						 "000111010010100110000000",
						 "000111010010100011001111",
						 "000111010010100000011110",
						 "000111010010011101101101",
						 "000111010010011010111100",
						 "000111010010011000001011",
						 "000111010010010101011010",
						 "000111010010010010101001",
						 "000111010010001111111000",
						 "000111010010001101000111",
						 "000111010010001010010110",
						 "000111010010000111100101",
						 "000111010010000100110100",
						 "000111010010000010000011",
						 "000111010001111111010010",
						 "000111010010101001000000",
						 "000111010010100110001110",
						 "000111010010100011011100",
						 "000111010010100000101010",
						 "000111010010011101111000",
						 "000111010010011011000110",
						 "000111010010011000010100",
						 "000111010010010101100010",
						 "000111010010010010110000",
						 "000111010010001111111110",
						 "000111010010001101001100",
						 "000111010010001010011010",
						 "000111010010000111101000",
						 "000111010010000100110110",
						 "000111010010000010000100",
						 "000111010001111111010010",
						 "000111010010101001000000",
						 "000111010010100110001110",
						 "000111010010100011011100",
						 "000111010010100000101010",
						 "000111010010011101111000",
						 "000111010010011011000110",
						 "000111010010011000010100",
						 "000111010010010101100010",
						 "000111010010010010110000",
						 "000111010010001111111110",
						 "000111010010001101001100",
						 "000111010010001010011010",
						 "000111010010000111101000",
						 "000111010010000100110110",
						 "000111010010000010000100",
						 "000111010001111111010010",
						 "000111010000000110000010",
						 "000111010000000011010000",
						 "000111010000000000011110",
						 "000111001111111101101100",
						 "000111001111111010111010",
						 "000111001111111000001000",
						 "000111001111110101010110",
						 "000111001111110010100100",
						 "000111001111101111110010",
						 "000111001111101101000000",
						 "000111001111101010001110",
						 "000111001111100111011100",
						 "000111001111100100101010",
						 "000111001111100001111000",
						 "000111001111011111000110",
						 "000111001111011100010100",
						 "000111010000000110010001",
						 "000111010000000011011110",
						 "000111010000000000101011",
						 "000111001111111101111000",
						 "000111001111111011000101",
						 "000111001111111000010010",
						 "000111001111110101011111",
						 "000111001111110010101100",
						 "000111001111101111111001",
						 "000111001111101101000110",
						 "000111001111101010010011",
						 "000111001111100111100000",
						 "000111001111100100101101",
						 "000111001111100001111010",
						 "000111001111011111000111",
						 "000111001111011100010100",
						 "000111010000000110010001",
						 "000111010000000011011110",
						 "000111010000000000101011",
						 "000111001111111101111000",
						 "000111001111111011000101",
						 "000111001111111000010010",
						 "000111001111110101011111",
						 "000111001111110010101100",
						 "000111001111101111111001",
						 "000111001111101101000110",
						 "000111001111101010010011",
						 "000111001111100111100000",
						 "000111001111100100101101",
						 "000111001111100001111010",
						 "000111001111011111000111",
						 "000111001111011100010100",
						 "000111001101100011010011",
						 "000111001101100000100000",
						 "000111001101011101101101",
						 "000111001101011010111010",
						 "000111001101011000000111",
						 "000111001101010101010100",
						 "000111001101010010100001",
						 "000111001101001111101110",
						 "000111001101001100111011",
						 "000111001101001010001000",
						 "000111001101000111010101",
						 "000111001101000100100010",
						 "000111001101000001101111",
						 "000111001100111110111100",
						 "000111001100111100001001",
						 "000111001100111001010110",
						 "000111001101100011010011",
						 "000111001101100000100000",
						 "000111001101011101101101",
						 "000111001101011010111010",
						 "000111001101011000000111",
						 "000111001101010101010100",
						 "000111001101010010100001",
						 "000111001101001111101110",
						 "000111001101001100111011",
						 "000111001101001010001000",
						 "000111001101000111010101",
						 "000111001101000100100010",
						 "000111001101000001101111",
						 "000111001100111110111100",
						 "000111001100111100001001",
						 "000111001100111001010110",
						 "000111001101100011100010",
						 "000111001101100000101110",
						 "000111001101011101111010",
						 "000111001101011011000110",
						 "000111001101011000010010",
						 "000111001101010101011110",
						 "000111001101010010101010",
						 "000111001101001111110110",
						 "000111001101001101000010",
						 "000111001101001010001110",
						 "000111001101000111011010",
						 "000111001101000100100110",
						 "000111001101000001110010",
						 "000111001100111110111110",
						 "000111001100111100001010",
						 "000111001100111001010110",
						 "000111001101100011100010",
						 "000111001101100000101110",
						 "000111001101011101111010",
						 "000111001101011011000110",
						 "000111001101011000010010",
						 "000111001101010101011110",
						 "000111001101010010101010",
						 "000111001101001111110110",
						 "000111001101001101000010",
						 "000111001101001010001110",
						 "000111001101000111011010",
						 "000111001101000100100110",
						 "000111001101000001110010",
						 "000111001100111110111110",
						 "000111001100111100001010",
						 "000111001100111001010110",
						 "000111001011000000100100",
						 "000111001010111101110000",
						 "000111001010111010111100",
						 "000111001010111000001000",
						 "000111001010110101010100",
						 "000111001010110010100000",
						 "000111001010101111101100",
						 "000111001010101100111000",
						 "000111001010101010000100",
						 "000111001010100111010000",
						 "000111001010100100011100",
						 "000111001010100001101000",
						 "000111001010011110110100",
						 "000111001010011100000000",
						 "000111001010011001001100",
						 "000111001010010110011000",
						 "000111001011000000100100",
						 "000111001010111101110000",
						 "000111001010111010111100",
						 "000111001010111000001000",
						 "000111001010110101010100",
						 "000111001010110010100000",
						 "000111001010101111101100",
						 "000111001010101100111000",
						 "000111001010101010000100",
						 "000111001010100111010000",
						 "000111001010100100011100",
						 "000111001010100001101000",
						 "000111001010011110110100",
						 "000111001010011100000000",
						 "000111001010011001001100",
						 "000111001010010110011000",
						 "000111001011000000110011",
						 "000111001010111101111110",
						 "000111001010111011001001",
						 "000111001010111000010100",
						 "000111001010110101011111",
						 "000111001010110010101010",
						 "000111001010101111110101",
						 "000111001010101101000000",
						 "000111001010101010001011",
						 "000111001010100111010110",
						 "000111001010100100100001",
						 "000111001010100001101100",
						 "000111001010011110110111",
						 "000111001010011100000010",
						 "000111001010011001001101",
						 "000111001010010110011000",
						 "000111001000011101110101",
						 "000111001000011011000000",
						 "000111001000011000001011",
						 "000111001000010101010110",
						 "000111001000010010100001",
						 "000111001000001111101100",
						 "000111001000001100110111",
						 "000111001000001010000010",
						 "000111001000000111001101",
						 "000111001000000100011000",
						 "000111001000000001100011",
						 "000111000111111110101110",
						 "000111000111111011111001",
						 "000111000111111001000100",
						 "000111000111110110001111",
						 "000111000111110011011010",
						 "000111001000011101110101",
						 "000111001000011011000000",
						 "000111001000011000001011",
						 "000111001000010101010110",
						 "000111001000010010100001",
						 "000111001000001111101100",
						 "000111001000001100110111",
						 "000111001000001010000010",
						 "000111001000000111001101",
						 "000111001000000100011000",
						 "000111001000000001100011",
						 "000111000111111110101110",
						 "000111000111111011111001",
						 "000111000111111001000100",
						 "000111000111110110001111",
						 "000111000111110011011010",
						 "000111001000011110000100",
						 "000111001000011011001110",
						 "000111001000011000011000",
						 "000111001000010101100010",
						 "000111001000010010101100",
						 "000111001000001111110110",
						 "000111001000001101000000",
						 "000111001000001010001010",
						 "000111001000000111010100",
						 "000111001000000100011110",
						 "000111001000000001101000",
						 "000111000111111110110010",
						 "000111000111111011111100",
						 "000111000111111001000110",
						 "000111000111110110010000",
						 "000111000111110011011010",
						 "000111001000011110000100",
						 "000111001000011011001110",
						 "000111001000011000011000",
						 "000111001000010101100010",
						 "000111001000010010101100",
						 "000111001000001111110110",
						 "000111001000001101000000",
						 "000111001000001010001010",
						 "000111001000000111010100",
						 "000111001000000100011110",
						 "000111001000000001101000",
						 "000111000111111110110010",
						 "000111000111111011111100",
						 "000111000111111001000110",
						 "000111000111110110010000",
						 "000111000111110011011010",
						 "000111000101111011000110",
						 "000111000101111000010000",
						 "000111000101110101011010",
						 "000111000101110010100100",
						 "000111000101101111101110",
						 "000111000101101100111000",
						 "000111000101101010000010",
						 "000111000101100111001100",
						 "000111000101100100010110",
						 "000111000101100001100000",
						 "000111000101011110101010",
						 "000111000101011011110100",
						 "000111000101011000111110",
						 "000111000101010110001000",
						 "000111000101010011010010",
						 "000111000101010000011100",
						 "000111000101111011000110",
						 "000111000101111000010000",
						 "000111000101110101011010",
						 "000111000101110010100100",
						 "000111000101101111101110",
						 "000111000101101100111000",
						 "000111000101101010000010",
						 "000111000101100111001100",
						 "000111000101100100010110",
						 "000111000101100001100000",
						 "000111000101011110101010",
						 "000111000101011011110100",
						 "000111000101011000111110",
						 "000111000101010110001000",
						 "000111000101010011010010",
						 "000111000101010000011100",
						 "000111000101111011010101",
						 "000111000101111000011110",
						 "000111000101110101100111",
						 "000111000101110010110000",
						 "000111000101101111111001",
						 "000111000101101101000010",
						 "000111000101101010001011",
						 "000111000101100111010100",
						 "000111000101100100011101",
						 "000111000101100001100110",
						 "000111000101011110101111",
						 "000111000101011011111000",
						 "000111000101011001000001",
						 "000111000101010110001010",
						 "000111000101010011010011",
						 "000111000101010000011100",
						 "000111000101111011010101",
						 "000111000101111000011110",
						 "000111000101110101100111",
						 "000111000101110010110000",
						 "000111000101101111111001",
						 "000111000101101101000010",
						 "000111000101101010001011",
						 "000111000101100111010100",
						 "000111000101100100011101",
						 "000111000101100001100110",
						 "000111000101011110101111",
						 "000111000101011011111000",
						 "000111000101011001000001",
						 "000111000101010110001010",
						 "000111000101010011010011",
						 "000111000101010000011100",
						 "000111000011011000010111",
						 "000111000011010101100000",
						 "000111000011010010101001",
						 "000111000011001111110010",
						 "000111000011001100111011",
						 "000111000011001010000100",
						 "000111000011000111001101",
						 "000111000011000100010110",
						 "000111000011000001011111",
						 "000111000010111110101000",
						 "000111000010111011110001",
						 "000111000010111000111010",
						 "000111000010110110000011",
						 "000111000010110011001100",
						 "000111000010110000010101",
						 "000111000010101101011110",
						 "000111000011011000010111",
						 "000111000011010101100000",
						 "000111000011010010101001",
						 "000111000011001111110010",
						 "000111000011001100111011",
						 "000111000011001010000100",
						 "000111000011000111001101",
						 "000111000011000100010110",
						 "000111000011000001011111",
						 "000111000010111110101000",
						 "000111000010111011110001",
						 "000111000010111000111010",
						 "000111000010110110000011",
						 "000111000010110011001100",
						 "000111000010110000010101",
						 "000111000010101101011110",
						 "000111000011011000100110",
						 "000111000011010101101110",
						 "000111000011010010110110",
						 "000111000011001111111110",
						 "000111000011001101000110",
						 "000111000011001010001110",
						 "000111000011000111010110",
						 "000111000011000100011110",
						 "000111000011000001100110",
						 "000111000010111110101110",
						 "000111000010111011110110",
						 "000111000010111000111110",
						 "000111000010110110000110",
						 "000111000010110011001110",
						 "000111000010110000010110",
						 "000111000010101101011110",
						 "000111000000110101101000",
						 "000111000000110010110000",
						 "000111000000101111111000",
						 "000111000000101101000000",
						 "000111000000101010001000",
						 "000111000000100111010000",
						 "000111000000100100011000",
						 "000111000000100001100000",
						 "000111000000011110101000",
						 "000111000000011011110000",
						 "000111000000011000111000",
						 "000111000000010110000000",
						 "000111000000010011001000",
						 "000111000000010000010000",
						 "000111000000001101011000",
						 "000111000000001010100000",
						 "000111000000110101101000",
						 "000111000000110010110000",
						 "000111000000101111111000",
						 "000111000000101101000000",
						 "000111000000101010001000",
						 "000111000000100111010000",
						 "000111000000100100011000",
						 "000111000000100001100000",
						 "000111000000011110101000",
						 "000111000000011011110000",
						 "000111000000011000111000",
						 "000111000000010110000000",
						 "000111000000010011001000",
						 "000111000000010000010000",
						 "000111000000001101011000",
						 "000111000000001010100000",
						 "000111000000110101110111",
						 "000111000000110010111110",
						 "000111000000110000000101",
						 "000111000000101101001100",
						 "000111000000101010010011",
						 "000111000000100111011010",
						 "000111000000100100100001",
						 "000111000000100001101000",
						 "000111000000011110101111",
						 "000111000000011011110110",
						 "000111000000011000111101",
						 "000111000000010110000100",
						 "000111000000010011001011",
						 "000111000000010000010010",
						 "000111000000001101011001",
						 "000111000000001010100000",
						 "000111000000110101110111",
						 "000111000000110010111110",
						 "000111000000110000000101",
						 "000111000000101101001100",
						 "000111000000101010010011",
						 "000111000000100111011010",
						 "000111000000100100100001",
						 "000111000000100001101000",
						 "000111000000011110101111",
						 "000111000000011011110110",
						 "000111000000011000111101",
						 "000111000000010110000100",
						 "000111000000010011001011",
						 "000111000000010000010010",
						 "000111000000001101011001",
						 "000111000000001010100000",
						 "000110111110010010111001",
						 "000110111110010000000000",
						 "000110111110001101000111",
						 "000110111110001010001110",
						 "000110111110000111010101",
						 "000110111110000100011100",
						 "000110111110000001100011",
						 "000110111101111110101010",
						 "000110111101111011110001",
						 "000110111101111000111000",
						 "000110111101110101111111",
						 "000110111101110011000110",
						 "000110111101110000001101",
						 "000110111101101101010100",
						 "000110111101101010011011",
						 "000110111101100111100010",
						 "000110111110010010111001",
						 "000110111110010000000000",
						 "000110111110001101000111",
						 "000110111110001010001110",
						 "000110111110000111010101",
						 "000110111110000100011100",
						 "000110111110000001100011",
						 "000110111101111110101010",
						 "000110111101111011110001",
						 "000110111101111000111000",
						 "000110111101110101111111",
						 "000110111101110011000110",
						 "000110111101110000001101",
						 "000110111101101101010100",
						 "000110111101101010011011",
						 "000110111101100111100010",
						 "000110111110010011001000",
						 "000110111110010000001110",
						 "000110111110001101010100",
						 "000110111110001010011010",
						 "000110111110000111100000",
						 "000110111110000100100110",
						 "000110111110000001101100",
						 "000110111101111110110010",
						 "000110111101111011111000",
						 "000110111101111000111110",
						 "000110111101110110000100",
						 "000110111101110011001010",
						 "000110111101110000010000",
						 "000110111101101101010110",
						 "000110111101101010011100",
						 "000110111101100111100010",
						 "000110111011110000001010",
						 "000110111011101101010000",
						 "000110111011101010010110",
						 "000110111011100111011100",
						 "000110111011100100100010",
						 "000110111011100001101000",
						 "000110111011011110101110",
						 "000110111011011011110100",
						 "000110111011011000111010",
						 "000110111011010110000000",
						 "000110111011010011000110",
						 "000110111011010000001100",
						 "000110111011001101010010",
						 "000110111011001010011000",
						 "000110111011000111011110",
						 "000110111011000100100100",
						 "000110111011110000001010",
						 "000110111011101101010000",
						 "000110111011101010010110",
						 "000110111011100111011100",
						 "000110111011100100100010",
						 "000110111011100001101000",
						 "000110111011011110101110",
						 "000110111011011011110100",
						 "000110111011011000111010",
						 "000110111011010110000000",
						 "000110111011010011000110",
						 "000110111011010000001100",
						 "000110111011001101010010",
						 "000110111011001010011000",
						 "000110111011000111011110",
						 "000110111011000100100100",
						 "000110111011110000001010",
						 "000110111011101101010000",
						 "000110111011101010010110",
						 "000110111011100111011100",
						 "000110111011100100100010",
						 "000110111011100001101000",
						 "000110111011011110101110",
						 "000110111011011011110100",
						 "000110111011011000111010",
						 "000110111011010110000000",
						 "000110111011010011000110",
						 "000110111011010000001100",
						 "000110111011001101010010",
						 "000110111011001010011000",
						 "000110111011000111011110",
						 "000110111011000100100100",
						 "000110111011110000011001",
						 "000110111011101101011110",
						 "000110111011101010100011",
						 "000110111011100111101000",
						 "000110111011100100101101",
						 "000110111011100001110010",
						 "000110111011011110110111",
						 "000110111011011011111100",
						 "000110111011011001000001",
						 "000110111011010110000110",
						 "000110111011010011001011",
						 "000110111011010000010000",
						 "000110111011001101010101",
						 "000110111011001010011010",
						 "000110111011000111011111",
						 "000110111011000100100100",
						 "000110111001001101011011",
						 "000110111001001010100000",
						 "000110111001000111100101",
						 "000110111001000100101010",
						 "000110111001000001101111",
						 "000110111000111110110100",
						 "000110111000111011111001",
						 "000110111000111000111110",
						 "000110111000110110000011",
						 "000110111000110011001000",
						 "000110111000110000001101",
						 "000110111000101101010010",
						 "000110111000101010010111",
						 "000110111000100111011100",
						 "000110111000100100100001",
						 "000110111000100001100110",
						 "000110111001001101011011",
						 "000110111001001010100000",
						 "000110111001000111100101",
						 "000110111001000100101010",
						 "000110111001000001101111",
						 "000110111000111110110100",
						 "000110111000111011111001",
						 "000110111000111000111110",
						 "000110111000110110000011",
						 "000110111000110011001000",
						 "000110111000110000001101",
						 "000110111000101101010010",
						 "000110111000101010010111",
						 "000110111000100111011100",
						 "000110111000100100100001",
						 "000110111000100001100110",
						 "000110111001001101011011",
						 "000110111001001010100000",
						 "000110111001000111100101",
						 "000110111001000100101010",
						 "000110111001000001101111",
						 "000110111000111110110100",
						 "000110111000111011111001",
						 "000110111000111000111110",
						 "000110111000110110000011",
						 "000110111000110011001000",
						 "000110111000110000001101",
						 "000110111000101101010010",
						 "000110111000101010010111",
						 "000110111000100111011100",
						 "000110111000100100100001",
						 "000110111000100001100110",
						 "000110110110101010101100",
						 "000110110110100111110000",
						 "000110110110100100110100",
						 "000110110110100001111000",
						 "000110110110011110111100",
						 "000110110110011100000000",
						 "000110110110011001000100",
						 "000110110110010110001000",
						 "000110110110010011001100",
						 "000110110110010000010000",
						 "000110110110001101010100",
						 "000110110110001010011000",
						 "000110110110000111011100",
						 "000110110110000100100000",
						 "000110110110000001100100",
						 "000110110101111110101000",
						 "000110110110101010101100",
						 "000110110110100111110000",
						 "000110110110100100110100",
						 "000110110110100001111000",
						 "000110110110011110111100",
						 "000110110110011100000000",
						 "000110110110011001000100",
						 "000110110110010110001000",
						 "000110110110010011001100",
						 "000110110110010000010000",
						 "000110110110001101010100",
						 "000110110110001010011000",
						 "000110110110000111011100",
						 "000110110110000100100000",
						 "000110110110000001100100",
						 "000110110101111110101000",
						 "000110110110101010101100",
						 "000110110110100111110000",
						 "000110110110100100110100",
						 "000110110110100001111000",
						 "000110110110011110111100",
						 "000110110110011100000000",
						 "000110110110011001000100",
						 "000110110110010110001000",
						 "000110110110010011001100",
						 "000110110110010000010000",
						 "000110110110001101010100",
						 "000110110110001010011000",
						 "000110110110000111011100",
						 "000110110110000100100000",
						 "000110110110000001100100",
						 "000110110101111110101000",
						 "000110110110101010111011",
						 "000110110110100111111110",
						 "000110110110100101000001",
						 "000110110110100010000100",
						 "000110110110011111000111",
						 "000110110110011100001010",
						 "000110110110011001001101",
						 "000110110110010110010000",
						 "000110110110010011010011",
						 "000110110110010000010110",
						 "000110110110001101011001",
						 "000110110110001010011100",
						 "000110110110000111011111",
						 "000110110110000100100010",
						 "000110110110000001100101",
						 "000110110101111110101000",
						 "000110110100000111111101",
						 "000110110100000101000000",
						 "000110110100000010000011",
						 "000110110011111111000110",
						 "000110110011111100001001",
						 "000110110011111001001100",
						 "000110110011110110001111",
						 "000110110011110011010010",
						 "000110110011110000010101",
						 "000110110011101101011000",
						 "000110110011101010011011",
						 "000110110011100111011110",
						 "000110110011100100100001",
						 "000110110011100001100100",
						 "000110110011011110100111",
						 "000110110011011011101010",
						 "000110110100000111111101",
						 "000110110100000101000000",
						 "000110110100000010000011",
						 "000110110011111111000110",
						 "000110110011111100001001",
						 "000110110011111001001100",
						 "000110110011110110001111",
						 "000110110011110011010010",
						 "000110110011110000010101",
						 "000110110011101101011000",
						 "000110110011101010011011",
						 "000110110011100111011110",
						 "000110110011100100100001",
						 "000110110011100001100100",
						 "000110110011011110100111",
						 "000110110011011011101010",
						 "000110110100000111111101",
						 "000110110100000101000000",
						 "000110110100000010000011",
						 "000110110011111111000110",
						 "000110110011111100001001",
						 "000110110011111001001100",
						 "000110110011110110001111",
						 "000110110011110011010010",
						 "000110110011110000010101",
						 "000110110011101101011000",
						 "000110110011101010011011",
						 "000110110011100111011110",
						 "000110110011100100100001",
						 "000110110011100001100100",
						 "000110110011011110100111",
						 "000110110011011011101010",
						 "000110110001100101001110",
						 "000110110001100010010000",
						 "000110110001011111010010",
						 "000110110001011100010100",
						 "000110110001011001010110",
						 "000110110001010110011000",
						 "000110110001010011011010",
						 "000110110001010000011100",
						 "000110110001001101011110",
						 "000110110001001010100000",
						 "000110110001000111100010",
						 "000110110001000100100100",
						 "000110110001000001100110",
						 "000110110000111110101000",
						 "000110110000111011101010",
						 "000110110000111000101100",
						 "000110110001100101001110",
						 "000110110001100010010000",
						 "000110110001011111010010",
						 "000110110001011100010100",
						 "000110110001011001010110",
						 "000110110001010110011000",
						 "000110110001010011011010",
						 "000110110001010000011100",
						 "000110110001001101011110",
						 "000110110001001010100000",
						 "000110110001000111100010",
						 "000110110001000100100100",
						 "000110110001000001100110",
						 "000110110000111110101000",
						 "000110110000111011101010",
						 "000110110000111000101100",
						 "000110110001100101001110",
						 "000110110001100010010000",
						 "000110110001011111010010",
						 "000110110001011100010100",
						 "000110110001011001010110",
						 "000110110001010110011000",
						 "000110110001010011011010",
						 "000110110001010000011100",
						 "000110110001001101011110",
						 "000110110001001010100000",
						 "000110110001000111100010",
						 "000110110001000100100100",
						 "000110110001000001100110",
						 "000110110000111110101000",
						 "000110110000111011101010",
						 "000110110000111000101100",
						 "000110110001100101001110",
						 "000110110001100010010000",
						 "000110110001011111010010",
						 "000110110001011100010100",
						 "000110110001011001010110",
						 "000110110001010110011000",
						 "000110110001010011011010",
						 "000110110001010000011100",
						 "000110110001001101011110",
						 "000110110001001010100000",
						 "000110110001000111100010",
						 "000110110001000100100100",
						 "000110110001000001100110",
						 "000110110000111110101000",
						 "000110110000111011101010",
						 "000110110000111000101100",
						 "000110101111000010011111",
						 "000110101110111111100000",
						 "000110101110111100100001",
						 "000110101110111001100010",
						 "000110101110110110100011",
						 "000110101110110011100100",
						 "000110101110110000100101",
						 "000110101110101101100110",
						 "000110101110101010100111",
						 "000110101110100111101000",
						 "000110101110100100101001",
						 "000110101110100001101010",
						 "000110101110011110101011",
						 "000110101110011011101100",
						 "000110101110011000101101",
						 "000110101110010101101110",
						 "000110101111000010011111",
						 "000110101110111111100000",
						 "000110101110111100100001",
						 "000110101110111001100010",
						 "000110101110110110100011",
						 "000110101110110011100100",
						 "000110101110110000100101",
						 "000110101110101101100110",
						 "000110101110101010100111",
						 "000110101110100111101000",
						 "000110101110100100101001",
						 "000110101110100001101010",
						 "000110101110011110101011",
						 "000110101110011011101100",
						 "000110101110011000101101",
						 "000110101110010101101110",
						 "000110101111000010011111",
						 "000110101110111111100000",
						 "000110101110111100100001",
						 "000110101110111001100010",
						 "000110101110110110100011",
						 "000110101110110011100100",
						 "000110101110110000100101",
						 "000110101110101101100110",
						 "000110101110101010100111",
						 "000110101110100111101000",
						 "000110101110100100101001",
						 "000110101110100001101010",
						 "000110101110011110101011",
						 "000110101110011011101100",
						 "000110101110011000101101",
						 "000110101110010101101110",
						 "000110101100011111100001",
						 "000110101100011100100010",
						 "000110101100011001100011",
						 "000110101100010110100100",
						 "000110101100010011100101",
						 "000110101100010000100110",
						 "000110101100001101100111",
						 "000110101100001010101000",
						 "000110101100000111101001",
						 "000110101100000100101010",
						 "000110101100000001101011",
						 "000110101011111110101100",
						 "000110101011111011101101",
						 "000110101011111000101110",
						 "000110101011110101101111",
						 "000110101011110010110000",
						 "000110101100011111110000",
						 "000110101100011100110000",
						 "000110101100011001110000",
						 "000110101100010110110000",
						 "000110101100010011110000",
						 "000110101100010000110000",
						 "000110101100001101110000",
						 "000110101100001010110000",
						 "000110101100000111110000",
						 "000110101100000100110000",
						 "000110101100000001110000",
						 "000110101011111110110000",
						 "000110101011111011110000",
						 "000110101011111000110000",
						 "000110101011110101110000",
						 "000110101011110010110000",
						 "000110101100011111110000",
						 "000110101100011100110000",
						 "000110101100011001110000",
						 "000110101100010110110000",
						 "000110101100010011110000",
						 "000110101100010000110000",
						 "000110101100001101110000",
						 "000110101100001010110000",
						 "000110101100000111110000",
						 "000110101100000100110000",
						 "000110101100000001110000",
						 "000110101011111110110000",
						 "000110101011111011110000",
						 "000110101011111000110000",
						 "000110101011110101110000",
						 "000110101011110010110000",
						 "000110101001111100110010",
						 "000110101001111001110010",
						 "000110101001110110110010",
						 "000110101001110011110010",
						 "000110101001110000110010",
						 "000110101001101101110010",
						 "000110101001101010110010",
						 "000110101001100111110010",
						 "000110101001100100110010",
						 "000110101001100001110010",
						 "000110101001011110110010",
						 "000110101001011011110010",
						 "000110101001011000110010",
						 "000110101001010101110010",
						 "000110101001010010110010",
						 "000110101001001111110010",
						 "000110101001111100110010",
						 "000110101001111001110010",
						 "000110101001110110110010",
						 "000110101001110011110010",
						 "000110101001110000110010",
						 "000110101001101101110010",
						 "000110101001101010110010",
						 "000110101001100111110010",
						 "000110101001100100110010",
						 "000110101001100001110010",
						 "000110101001011110110010",
						 "000110101001011011110010",
						 "000110101001011000110010",
						 "000110101001010101110010",
						 "000110101001010010110010",
						 "000110101001001111110010",
						 "000110101001111101000001",
						 "000110101001111010000000",
						 "000110101001110110111111",
						 "000110101001110011111110",
						 "000110101001110000111101",
						 "000110101001101101111100",
						 "000110101001101010111011",
						 "000110101001100111111010",
						 "000110101001100100111001",
						 "000110101001100001111000",
						 "000110101001011110110111",
						 "000110101001011011110110",
						 "000110101001011000110101",
						 "000110101001010101110100",
						 "000110101001010010110011",
						 "000110101001001111110010",
						 "000110101001111101000001",
						 "000110101001111010000000",
						 "000110101001110110111111",
						 "000110101001110011111110",
						 "000110101001110000111101",
						 "000110101001101101111100",
						 "000110101001101010111011",
						 "000110101001100111111010",
						 "000110101001100100111001",
						 "000110101001100001111000",
						 "000110101001011110110111",
						 "000110101001011011110110",
						 "000110101001011000110101",
						 "000110101001010101110100",
						 "000110101001010010110011",
						 "000110101001001111110010",
						 "000110100111011010000011",
						 "000110100111010111000010",
						 "000110100111010100000001",
						 "000110100111010001000000",
						 "000110100111001101111111",
						 "000110100111001010111110",
						 "000110100111000111111101",
						 "000110100111000100111100",
						 "000110100111000001111011",
						 "000110100110111110111010",
						 "000110100110111011111001",
						 "000110100110111000111000",
						 "000110100110110101110111",
						 "000110100110110010110110",
						 "000110100110101111110101",
						 "000110100110101100110100",
						 "000110100111011010000011",
						 "000110100111010111000010",
						 "000110100111010100000001",
						 "000110100111010001000000",
						 "000110100111001101111111",
						 "000110100111001010111110",
						 "000110100111000111111101",
						 "000110100111000100111100",
						 "000110100111000001111011",
						 "000110100110111110111010",
						 "000110100110111011111001",
						 "000110100110111000111000",
						 "000110100110110101110111",
						 "000110100110110010110110",
						 "000110100110101111110101",
						 "000110100110101100110100",
						 "000110100111011010010010",
						 "000110100111010111010000",
						 "000110100111010100001110",
						 "000110100111010001001100",
						 "000110100111001110001010",
						 "000110100111001011001000",
						 "000110100111001000000110",
						 "000110100111000101000100",
						 "000110100111000010000010",
						 "000110100110111111000000",
						 "000110100110111011111110",
						 "000110100110111000111100",
						 "000110100110110101111010",
						 "000110100110110010111000",
						 "000110100110101111110110",
						 "000110100110101100110100",
						 "000110100100110111010100",
						 "000110100100110100010010",
						 "000110100100110001010000",
						 "000110100100101110001110",
						 "000110100100101011001100",
						 "000110100100101000001010",
						 "000110100100100101001000",
						 "000110100100100010000110",
						 "000110100100011111000100",
						 "000110100100011100000010",
						 "000110100100011001000000",
						 "000110100100010101111110",
						 "000110100100010010111100",
						 "000110100100001111111010",
						 "000110100100001100111000",
						 "000110100100001001110110",
						 "000110100100110111010100",
						 "000110100100110100010010",
						 "000110100100110001010000",
						 "000110100100101110001110",
						 "000110100100101011001100",
						 "000110100100101000001010",
						 "000110100100100101001000",
						 "000110100100100010000110",
						 "000110100100011111000100",
						 "000110100100011100000010",
						 "000110100100011001000000",
						 "000110100100010101111110",
						 "000110100100010010111100",
						 "000110100100001111111010",
						 "000110100100001100111000",
						 "000110100100001001110110",
						 "000110100100110111010100",
						 "000110100100110100010010",
						 "000110100100110001010000",
						 "000110100100101110001110",
						 "000110100100101011001100",
						 "000110100100101000001010",
						 "000110100100100101001000",
						 "000110100100100010000110",
						 "000110100100011111000100",
						 "000110100100011100000010",
						 "000110100100011001000000",
						 "000110100100010101111110",
						 "000110100100010010111100",
						 "000110100100001111111010",
						 "000110100100001100111000",
						 "000110100100001001110110",
						 "000110100010010100100101",
						 "000110100010010001100010",
						 "000110100010001110011111",
						 "000110100010001011011100",
						 "000110100010001000011001",
						 "000110100010000101010110",
						 "000110100010000010010011",
						 "000110100001111111010000",
						 "000110100001111100001101",
						 "000110100001111001001010",
						 "000110100001110110000111",
						 "000110100001110011000100",
						 "000110100001110000000001",
						 "000110100001101100111110",
						 "000110100001101001111011",
						 "000110100001100110111000",
						 "000110100010010100100101",
						 "000110100010010001100010",
						 "000110100010001110011111",
						 "000110100010001011011100",
						 "000110100010001000011001",
						 "000110100010000101010110",
						 "000110100010000010010011",
						 "000110100001111111010000",
						 "000110100001111100001101",
						 "000110100001111001001010",
						 "000110100001110110000111",
						 "000110100001110011000100",
						 "000110100001110000000001",
						 "000110100001101100111110",
						 "000110100001101001111011",
						 "000110100001100110111000",
						 "000110100010010100100101",
						 "000110100010010001100010",
						 "000110100010001110011111",
						 "000110100010001011011100",
						 "000110100010001000011001",
						 "000110100010000101010110",
						 "000110100010000010010011",
						 "000110100001111111010000",
						 "000110100001111100001101",
						 "000110100001111001001010",
						 "000110100001110110000111",
						 "000110100001110011000100",
						 "000110100001110000000001",
						 "000110100001101100111110",
						 "000110100001101001111011",
						 "000110100001100110111000",
						 "000110100010010100100101",
						 "000110100010010001100010",
						 "000110100010001110011111",
						 "000110100010001011011100",
						 "000110100010001000011001",
						 "000110100010000101010110",
						 "000110100010000010010011",
						 "000110100001111111010000",
						 "000110100001111100001101",
						 "000110100001111001001010",
						 "000110100001110110000111",
						 "000110100001110011000100",
						 "000110100001110000000001",
						 "000110100001101100111110",
						 "000110100001101001111011",
						 "000110100001100110111000",
						 "000110011111110001110110",
						 "000110011111101110110010",
						 "000110011111101011101110",
						 "000110011111101000101010",
						 "000110011111100101100110",
						 "000110011111100010100010",
						 "000110011111011111011110",
						 "000110011111011100011010",
						 "000110011111011001010110",
						 "000110011111010110010010",
						 "000110011111010011001110",
						 "000110011111010000001010",
						 "000110011111001101000110",
						 "000110011111001010000010",
						 "000110011111000110111110",
						 "000110011111000011111010",
						 "000110011111110001110110",
						 "000110011111101110110010",
						 "000110011111101011101110",
						 "000110011111101000101010",
						 "000110011111100101100110",
						 "000110011111100010100010",
						 "000110011111011111011110",
						 "000110011111011100011010",
						 "000110011111011001010110",
						 "000110011111010110010010",
						 "000110011111010011001110",
						 "000110011111010000001010",
						 "000110011111001101000110",
						 "000110011111001010000010",
						 "000110011111000110111110",
						 "000110011111000011111010",
						 "000110011111110001110110",
						 "000110011111101110110010",
						 "000110011111101011101110",
						 "000110011111101000101010",
						 "000110011111100101100110",
						 "000110011111100010100010",
						 "000110011111011111011110",
						 "000110011111011100011010",
						 "000110011111011001010110",
						 "000110011111010110010010",
						 "000110011111010011001110",
						 "000110011111010000001010",
						 "000110011111001101000110",
						 "000110011111001010000010",
						 "000110011111000110111110",
						 "000110011111000011111010",
						 "000110011101001110111000",
						 "000110011101001011110100",
						 "000110011101001000110000",
						 "000110011101000101101100",
						 "000110011101000010101000",
						 "000110011100111111100100",
						 "000110011100111100100000",
						 "000110011100111001011100",
						 "000110011100110110011000",
						 "000110011100110011010100",
						 "000110011100110000010000",
						 "000110011100101101001100",
						 "000110011100101010001000",
						 "000110011100100111000100",
						 "000110011100100100000000",
						 "000110011100100000111100",
						 "000110011101001111000111",
						 "000110011101001100000010",
						 "000110011101001000111101",
						 "000110011101000101111000",
						 "000110011101000010110011",
						 "000110011100111111101110",
						 "000110011100111100101001",
						 "000110011100111001100100",
						 "000110011100110110011111",
						 "000110011100110011011010",
						 "000110011100110000010101",
						 "000110011100101101010000",
						 "000110011100101010001011",
						 "000110011100100111000110",
						 "000110011100100100000001",
						 "000110011100100000111100",
						 "000110011101001111000111",
						 "000110011101001100000010",
						 "000110011101001000111101",
						 "000110011101000101111000",
						 "000110011101000010110011",
						 "000110011100111111101110",
						 "000110011100111100101001",
						 "000110011100111001100100",
						 "000110011100110110011111",
						 "000110011100110011011010",
						 "000110011100110000010101",
						 "000110011100101101010000",
						 "000110011100101010001011",
						 "000110011100100111000110",
						 "000110011100100100000001",
						 "000110011100100000111100",
						 "000110011010101100001001",
						 "000110011010101001000100",
						 "000110011010100101111111",
						 "000110011010100010111010",
						 "000110011010011111110101",
						 "000110011010011100110000",
						 "000110011010011001101011",
						 "000110011010010110100110",
						 "000110011010010011100001",
						 "000110011010010000011100",
						 "000110011010001101010111",
						 "000110011010001010010010",
						 "000110011010000111001101",
						 "000110011010000100001000",
						 "000110011010000001000011",
						 "000110011001111101111110",
						 "000110011010101100001001",
						 "000110011010101001000100",
						 "000110011010100101111111",
						 "000110011010100010111010",
						 "000110011010011111110101",
						 "000110011010011100110000",
						 "000110011010011001101011",
						 "000110011010010110100110",
						 "000110011010010011100001",
						 "000110011010010000011100",
						 "000110011010001101010111",
						 "000110011010001010010010",
						 "000110011010000111001101",
						 "000110011010000100001000",
						 "000110011010000001000011",
						 "000110011001111101111110",
						 "000110011010101100011000",
						 "000110011010101001010010",
						 "000110011010100110001100",
						 "000110011010100011000110",
						 "000110011010100000000000",
						 "000110011010011100111010",
						 "000110011010011001110100",
						 "000110011010010110101110",
						 "000110011010010011101000",
						 "000110011010010000100010",
						 "000110011010001101011100",
						 "000110011010001010010110",
						 "000110011010000111010000",
						 "000110011010000100001010",
						 "000110011010000001000100",
						 "000110011001111101111110",
						 "000110011010101100011000",
						 "000110011010101001010010",
						 "000110011010100110001100",
						 "000110011010100011000110",
						 "000110011010100000000000",
						 "000110011010011100111010",
						 "000110011010011001110100",
						 "000110011010010110101110",
						 "000110011010010011101000",
						 "000110011010010000100010",
						 "000110011010001101011100",
						 "000110011010001010010110",
						 "000110011010000111010000",
						 "000110011010000100001010",
						 "000110011010000001000100",
						 "000110011001111101111110",
						 "000110011000001001011010",
						 "000110011000000110010100",
						 "000110011000000011001110",
						 "000110011000000000001000",
						 "000110010111111101000010",
						 "000110010111111001111100",
						 "000110010111110110110110",
						 "000110010111110011110000",
						 "000110010111110000101010",
						 "000110010111101101100100",
						 "000110010111101010011110",
						 "000110010111100111011000",
						 "000110010111100100010010",
						 "000110010111100001001100",
						 "000110010111011110000110",
						 "000110010111011011000000",
						 "000110011000001001011010",
						 "000110011000000110010100",
						 "000110011000000011001110",
						 "000110011000000000001000",
						 "000110010111111101000010",
						 "000110010111111001111100",
						 "000110010111110110110110",
						 "000110010111110011110000",
						 "000110010111110000101010",
						 "000110010111101101100100",
						 "000110010111101010011110",
						 "000110010111100111011000",
						 "000110010111100100010010",
						 "000110010111100001001100",
						 "000110010111011110000110",
						 "000110010111011011000000",
						 "000110011000001001101001",
						 "000110011000000110100010",
						 "000110011000000011011011",
						 "000110011000000000010100",
						 "000110010111111101001101",
						 "000110010111111010000110",
						 "000110010111110110111111",
						 "000110010111110011111000",
						 "000110010111110000110001",
						 "000110010111101101101010",
						 "000110010111101010100011",
						 "000110010111100111011100",
						 "000110010111100100010101",
						 "000110010111100001001110",
						 "000110010111011110000111",
						 "000110010111011011000000",
						 "000110010101100110101011",
						 "000110010101100011100100",
						 "000110010101100000011101",
						 "000110010101011101010110",
						 "000110010101011010001111",
						 "000110010101010111001000",
						 "000110010101010100000001",
						 "000110010101010000111010",
						 "000110010101001101110011",
						 "000110010101001010101100",
						 "000110010101000111100101",
						 "000110010101000100011110",
						 "000110010101000001010111",
						 "000110010100111110010000",
						 "000110010100111011001001",
						 "000110010100111000000010",
						 "000110010101100110101011",
						 "000110010101100011100100",
						 "000110010101100000011101",
						 "000110010101011101010110",
						 "000110010101011010001111",
						 "000110010101010111001000",
						 "000110010101010100000001",
						 "000110010101010000111010",
						 "000110010101001101110011",
						 "000110010101001010101100",
						 "000110010101000111100101",
						 "000110010101000100011110",
						 "000110010101000001010111",
						 "000110010100111110010000",
						 "000110010100111011001001",
						 "000110010100111000000010",
						 "000110010101100110101011",
						 "000110010101100011100100",
						 "000110010101100000011101",
						 "000110010101011101010110",
						 "000110010101011010001111",
						 "000110010101010111001000",
						 "000110010101010100000001",
						 "000110010101010000111010",
						 "000110010101001101110011",
						 "000110010101001010101100",
						 "000110010101000111100101",
						 "000110010101000100011110",
						 "000110010101000001010111",
						 "000110010100111110010000",
						 "000110010100111011001001",
						 "000110010100111000000010",
						 "000110010011000011111100",
						 "000110010011000000110100",
						 "000110010010111101101100",
						 "000110010010111010100100",
						 "000110010010110111011100",
						 "000110010010110100010100",
						 "000110010010110001001100",
						 "000110010010101110000100",
						 "000110010010101010111100",
						 "000110010010100111110100",
						 "000110010010100100101100",
						 "000110010010100001100100",
						 "000110010010011110011100",
						 "000110010010011011010100",
						 "000110010010011000001100",
						 "000110010010010101000100",
						 "000110010011000011111100",
						 "000110010011000000110100",
						 "000110010010111101101100",
						 "000110010010111010100100",
						 "000110010010110111011100",
						 "000110010010110100010100",
						 "000110010010110001001100",
						 "000110010010101110000100",
						 "000110010010101010111100",
						 "000110010010100111110100",
						 "000110010010100100101100",
						 "000110010010100001100100",
						 "000110010010011110011100",
						 "000110010010011011010100",
						 "000110010010011000001100",
						 "000110010010010101000100",
						 "000110010011000011111100",
						 "000110010011000000110100",
						 "000110010010111101101100",
						 "000110010010111010100100",
						 "000110010010110111011100",
						 "000110010010110100010100",
						 "000110010010110001001100",
						 "000110010010101110000100",
						 "000110010010101010111100",
						 "000110010010100111110100",
						 "000110010010100100101100",
						 "000110010010100001100100",
						 "000110010010011110011100",
						 "000110010010011011010100",
						 "000110010010011000001100",
						 "000110010010010101000100",
						 "000110010011000011111100",
						 "000110010011000000110100",
						 "000110010010111101101100",
						 "000110010010111010100100",
						 "000110010010110111011100",
						 "000110010010110100010100",
						 "000110010010110001001100",
						 "000110010010101110000100",
						 "000110010010101010111100",
						 "000110010010100111110100",
						 "000110010010100100101100",
						 "000110010010100001100100",
						 "000110010010011110011100",
						 "000110010010011011010100",
						 "000110010010011000001100",
						 "000110010010010101000100",
						 "000110010000100001001101",
						 "000110010000011110000100",
						 "000110010000011010111011",
						 "000110010000010111110010",
						 "000110010000010100101001",
						 "000110010000010001100000",
						 "000110010000001110010111",
						 "000110010000001011001110",
						 "000110010000001000000101",
						 "000110010000000100111100",
						 "000110010000000001110011",
						 "000110001111111110101010",
						 "000110001111111011100001",
						 "000110001111111000011000",
						 "000110001111110101001111",
						 "000110001111110010000110",
						 "000110010000100001001101",
						 "000110010000011110000100",
						 "000110010000011010111011",
						 "000110010000010111110010",
						 "000110010000010100101001",
						 "000110010000010001100000",
						 "000110010000001110010111",
						 "000110010000001011001110",
						 "000110010000001000000101",
						 "000110010000000100111100",
						 "000110010000000001110011",
						 "000110001111111110101010",
						 "000110001111111011100001",
						 "000110001111111000011000",
						 "000110001111110101001111",
						 "000110001111110010000110",
						 "000110010000100001001101",
						 "000110010000011110000100",
						 "000110010000011010111011",
						 "000110010000010111110010",
						 "000110010000010100101001",
						 "000110010000010001100000",
						 "000110010000001110010111",
						 "000110010000001011001110",
						 "000110010000001000000101",
						 "000110010000000100111100",
						 "000110010000000001110011",
						 "000110001111111110101010",
						 "000110001111111011100001",
						 "000110001111111000011000",
						 "000110001111110101001111",
						 "000110001111110010000110",
						 "000110001101111110001111",
						 "000110001101111011000110",
						 "000110001101110111111101",
						 "000110001101110100110100",
						 "000110001101110001101011",
						 "000110001101101110100010",
						 "000110001101101011011001",
						 "000110001101101000010000",
						 "000110001101100101000111",
						 "000110001101100001111110",
						 "000110001101011110110101",
						 "000110001101011011101100",
						 "000110001101011000100011",
						 "000110001101010101011010",
						 "000110001101010010010001",
						 "000110001101001111001000",
						 "000110001101111110011110",
						 "000110001101111011010100",
						 "000110001101111000001010",
						 "000110001101110101000000",
						 "000110001101110001110110",
						 "000110001101101110101100",
						 "000110001101101011100010",
						 "000110001101101000011000",
						 "000110001101100101001110",
						 "000110001101100010000100",
						 "000110001101011110111010",
						 "000110001101011011110000",
						 "000110001101011000100110",
						 "000110001101010101011100",
						 "000110001101010010010010",
						 "000110001101001111001000",
						 "000110001101111110011110",
						 "000110001101111011010100",
						 "000110001101111000001010",
						 "000110001101110101000000",
						 "000110001101110001110110",
						 "000110001101101110101100",
						 "000110001101101011100010",
						 "000110001101101000011000",
						 "000110001101100101001110",
						 "000110001101100010000100",
						 "000110001101011110111010",
						 "000110001101011011110000",
						 "000110001101011000100110",
						 "000110001101010101011100",
						 "000110001101010010010010",
						 "000110001101001111001000",
						 "000110001011011011100000",
						 "000110001011011000010110",
						 "000110001011010101001100",
						 "000110001011010010000010",
						 "000110001011001110111000",
						 "000110001011001011101110",
						 "000110001011001000100100",
						 "000110001011000101011010",
						 "000110001011000010010000",
						 "000110001010111111000110",
						 "000110001010111011111100",
						 "000110001010111000110010",
						 "000110001010110101101000",
						 "000110001010110010011110",
						 "000110001010101111010100",
						 "000110001010101100001010",
						 "000110001011011011100000",
						 "000110001011011000010110",
						 "000110001011010101001100",
						 "000110001011010010000010",
						 "000110001011001110111000",
						 "000110001011001011101110",
						 "000110001011001000100100",
						 "000110001011000101011010",
						 "000110001011000010010000",
						 "000110001010111111000110",
						 "000110001010111011111100",
						 "000110001010111000110010",
						 "000110001010110101101000",
						 "000110001010110010011110",
						 "000110001010101111010100",
						 "000110001010101100001010",
						 "000110001011011011101111",
						 "000110001011011000100100",
						 "000110001011010101011001",
						 "000110001011010010001110",
						 "000110001011001111000011",
						 "000110001011001011111000",
						 "000110001011001000101101",
						 "000110001011000101100010",
						 "000110001011000010010111",
						 "000110001010111111001100",
						 "000110001010111100000001",
						 "000110001010111000110110",
						 "000110001010110101101011",
						 "000110001010110010100000",
						 "000110001010101111010101",
						 "000110001010101100001010",
						 "000110001000111000110001",
						 "000110001000110101100110",
						 "000110001000110010011011",
						 "000110001000101111010000",
						 "000110001000101100000101",
						 "000110001000101000111010",
						 "000110001000100101101111",
						 "000110001000100010100100",
						 "000110001000011111011001",
						 "000110001000011100001110",
						 "000110001000011001000011",
						 "000110001000010101111000",
						 "000110001000010010101101",
						 "000110001000001111100010",
						 "000110001000001100010111",
						 "000110001000001001001100",
						 "000110001000111000110001",
						 "000110001000110101100110",
						 "000110001000110010011011",
						 "000110001000101111010000",
						 "000110001000101100000101",
						 "000110001000101000111010",
						 "000110001000100101101111",
						 "000110001000100010100100",
						 "000110001000011111011001",
						 "000110001000011100001110",
						 "000110001000011001000011",
						 "000110001000010101111000",
						 "000110001000010010101101",
						 "000110001000001111100010",
						 "000110001000001100010111",
						 "000110001000001001001100",
						 "000110001000111000110001",
						 "000110001000110101100110",
						 "000110001000110010011011",
						 "000110001000101111010000",
						 "000110001000101100000101",
						 "000110001000101000111010",
						 "000110001000100101101111",
						 "000110001000100010100100",
						 "000110001000011111011001",
						 "000110001000011100001110",
						 "000110001000011001000011",
						 "000110001000010101111000",
						 "000110001000010010101101",
						 "000110001000001111100010",
						 "000110001000001100010111",
						 "000110001000001001001100",
						 "000110000110010110000010",
						 "000110000110010010110110",
						 "000110000110001111101010",
						 "000110000110001100011110",
						 "000110000110001001010010",
						 "000110000110000110000110",
						 "000110000110000010111010",
						 "000110000101111111101110",
						 "000110000101111100100010",
						 "000110000101111001010110",
						 "000110000101110110001010",
						 "000110000101110010111110",
						 "000110000101101111110010",
						 "000110000101101100100110",
						 "000110000101101001011010",
						 "000110000101100110001110",
						 "000110000110010110000010",
						 "000110000110010010110110",
						 "000110000110001111101010",
						 "000110000110001100011110",
						 "000110000110001001010010",
						 "000110000110000110000110",
						 "000110000110000010111010",
						 "000110000101111111101110",
						 "000110000101111100100010",
						 "000110000101111001010110",
						 "000110000101110110001010",
						 "000110000101110010111110",
						 "000110000101101111110010",
						 "000110000101101100100110",
						 "000110000101101001011010",
						 "000110000101100110001110",
						 "000110000110010110000010",
						 "000110000110010010110110",
						 "000110000110001111101010",
						 "000110000110001100011110",
						 "000110000110001001010010",
						 "000110000110000110000110",
						 "000110000110000010111010",
						 "000110000101111111101110",
						 "000110000101111100100010",
						 "000110000101111001010110",
						 "000110000101110110001010",
						 "000110000101110010111110",
						 "000110000101101111110010",
						 "000110000101101100100110",
						 "000110000101101001011010",
						 "000110000101100110001110",
						 "000110000110010110000010",
						 "000110000110010010110110",
						 "000110000110001111101010",
						 "000110000110001100011110",
						 "000110000110001001010010",
						 "000110000110000110000110",
						 "000110000110000010111010",
						 "000110000101111111101110",
						 "000110000101111100100010",
						 "000110000101111001010110",
						 "000110000101110110001010",
						 "000110000101110010111110",
						 "000110000101101111110010",
						 "000110000101101100100110",
						 "000110000101101001011010",
						 "000110000101100110001110",
						 "000110000011110011000100",
						 "000110000011101111111000",
						 "000110000011101100101100",
						 "000110000011101001100000",
						 "000110000011100110010100",
						 "000110000011100011001000",
						 "000110000011011111111100",
						 "000110000011011100110000",
						 "000110000011011001100100",
						 "000110000011010110011000",
						 "000110000011010011001100",
						 "000110000011010000000000",
						 "000110000011001100110100",
						 "000110000011001001101000",
						 "000110000011000110011100",
						 "000110000011000011010000",
						 "000110000011110011010011",
						 "000110000011110000000110",
						 "000110000011101100111001",
						 "000110000011101001101100",
						 "000110000011100110011111",
						 "000110000011100011010010",
						 "000110000011100000000101",
						 "000110000011011100111000",
						 "000110000011011001101011",
						 "000110000011010110011110",
						 "000110000011010011010001",
						 "000110000011010000000100",
						 "000110000011001100110111",
						 "000110000011001001101010",
						 "000110000011000110011101",
						 "000110000011000011010000",
						 "000110000011110011010011",
						 "000110000011110000000110",
						 "000110000011101100111001",
						 "000110000011101001101100",
						 "000110000011100110011111",
						 "000110000011100011010010",
						 "000110000011100000000101",
						 "000110000011011100111000",
						 "000110000011011001101011",
						 "000110000011010110011110",
						 "000110000011010011010001",
						 "000110000011010000000100",
						 "000110000011001100110111",
						 "000110000011001001101010",
						 "000110000011000110011101",
						 "000110000011000011010000",
						 "000110000001010000010101",
						 "000110000001001101001000",
						 "000110000001001001111011",
						 "000110000001000110101110",
						 "000110000001000011100001",
						 "000110000001000000010100",
						 "000110000000111101000111",
						 "000110000000111001111010",
						 "000110000000110110101101",
						 "000110000000110011100000",
						 "000110000000110000010011",
						 "000110000000101101000110",
						 "000110000000101001111001",
						 "000110000000100110101100",
						 "000110000000100011011111",
						 "000110000000100000010010",
						 "000110000001010000010101",
						 "000110000001001101001000",
						 "000110000001001001111011",
						 "000110000001000110101110",
						 "000110000001000011100001",
						 "000110000001000000010100",
						 "000110000000111101000111",
						 "000110000000111001111010",
						 "000110000000110110101101",
						 "000110000000110011100000",
						 "000110000000110000010011",
						 "000110000000101101000110",
						 "000110000000101001111001",
						 "000110000000100110101100",
						 "000110000000100011011111",
						 "000110000000100000010010",
						 "000110000001010000100100",
						 "000110000001001101010110",
						 "000110000001001010001000",
						 "000110000001000110111010",
						 "000110000001000011101100",
						 "000110000001000000011110",
						 "000110000000111101010000",
						 "000110000000111010000010",
						 "000110000000110110110100",
						 "000110000000110011100110",
						 "000110000000110000011000",
						 "000110000000101101001010",
						 "000110000000101001111100",
						 "000110000000100110101110",
						 "000110000000100011100000",
						 "000110000000100000010010",
						 "000101111110101101100110",
						 "000101111110101010011000",
						 "000101111110100111001010",
						 "000101111110100011111100",
						 "000101111110100000101110",
						 "000101111110011101100000",
						 "000101111110011010010010",
						 "000101111110010111000100",
						 "000101111110010011110110",
						 "000101111110010000101000",
						 "000101111110001101011010",
						 "000101111110001010001100",
						 "000101111110000110111110",
						 "000101111110000011110000",
						 "000101111110000000100010",
						 "000101111101111101010100",
						 "000101111110101101100110",
						 "000101111110101010011000",
						 "000101111110100111001010",
						 "000101111110100011111100",
						 "000101111110100000101110",
						 "000101111110011101100000",
						 "000101111110011010010010",
						 "000101111110010111000100",
						 "000101111110010011110110",
						 "000101111110010000101000",
						 "000101111110001101011010",
						 "000101111110001010001100",
						 "000101111110000110111110",
						 "000101111110000011110000",
						 "000101111110000000100010",
						 "000101111101111101010100",
						 "000101111110101101100110",
						 "000101111110101010011000",
						 "000101111110100111001010",
						 "000101111110100011111100",
						 "000101111110100000101110",
						 "000101111110011101100000",
						 "000101111110011010010010",
						 "000101111110010111000100",
						 "000101111110010011110110",
						 "000101111110010000101000",
						 "000101111110001101011010",
						 "000101111110001010001100",
						 "000101111110000110111110",
						 "000101111110000011110000",
						 "000101111110000000100010",
						 "000101111101111101010100",
						 "000101111100001010110111",
						 "000101111100000111101000",
						 "000101111100000100011001",
						 "000101111100000001001010",
						 "000101111011111101111011",
						 "000101111011111010101100",
						 "000101111011110111011101",
						 "000101111011110100001110",
						 "000101111011110000111111",
						 "000101111011101101110000",
						 "000101111011101010100001",
						 "000101111011100111010010",
						 "000101111011100100000011",
						 "000101111011100000110100",
						 "000101111011011101100101",
						 "000101111011011010010110",
						 "000101111100001010110111",
						 "000101111100000111101000",
						 "000101111100000100011001",
						 "000101111100000001001010",
						 "000101111011111101111011",
						 "000101111011111010101100",
						 "000101111011110111011101",
						 "000101111011110100001110",
						 "000101111011110000111111",
						 "000101111011101101110000",
						 "000101111011101010100001",
						 "000101111011100111010010",
						 "000101111011100100000011",
						 "000101111011100000110100",
						 "000101111011011101100101",
						 "000101111011011010010110",
						 "000101111100001010110111",
						 "000101111100000111101000",
						 "000101111100000100011001",
						 "000101111100000001001010",
						 "000101111011111101111011",
						 "000101111011111010101100",
						 "000101111011110111011101",
						 "000101111011110100001110",
						 "000101111011110000111111",
						 "000101111011101101110000",
						 "000101111011101010100001",
						 "000101111011100111010010",
						 "000101111011100100000011",
						 "000101111011100000110100",
						 "000101111011011101100101",
						 "000101111011011010010110",
						 "000101111001100111111001",
						 "000101111001100100101010",
						 "000101111001100001011011",
						 "000101111001011110001100",
						 "000101111001011010111101",
						 "000101111001010111101110",
						 "000101111001010100011111",
						 "000101111001010001010000",
						 "000101111001001110000001",
						 "000101111001001010110010",
						 "000101111001000111100011",
						 "000101111001000100010100",
						 "000101111001000001000101",
						 "000101111000111101110110",
						 "000101111000111010100111",
						 "000101111000110111011000",
						 "000101111001100111111001",
						 "000101111001100100101010",
						 "000101111001100001011011",
						 "000101111001011110001100",
						 "000101111001011010111101",
						 "000101111001010111101110",
						 "000101111001010100011111",
						 "000101111001010001010000",
						 "000101111001001110000001",
						 "000101111001001010110010",
						 "000101111001000111100011",
						 "000101111001000100010100",
						 "000101111001000001000101",
						 "000101111000111101110110",
						 "000101111000111010100111",
						 "000101111000110111011000",
						 "000101111001101000001000",
						 "000101111001100100111000",
						 "000101111001100001101000",
						 "000101111001011110011000",
						 "000101111001011011001000",
						 "000101111001010111111000",
						 "000101111001010100101000",
						 "000101111001010001011000",
						 "000101111001001110001000",
						 "000101111001001010111000",
						 "000101111001000111101000",
						 "000101111001000100011000",
						 "000101111001000001001000",
						 "000101111000111101111000",
						 "000101111000111010101000",
						 "000101111000110111011000",
						 "000101110111000101001010",
						 "000101110111000001111010",
						 "000101110110111110101010",
						 "000101110110111011011010",
						 "000101110110111000001010",
						 "000101110110110100111010",
						 "000101110110110001101010",
						 "000101110110101110011010",
						 "000101110110101011001010",
						 "000101110110100111111010",
						 "000101110110100100101010",
						 "000101110110100001011010",
						 "000101110110011110001010",
						 "000101110110011010111010",
						 "000101110110010111101010",
						 "000101110110010100011010",
						 "000101110111000101001010",
						 "000101110111000001111010",
						 "000101110110111110101010",
						 "000101110110111011011010",
						 "000101110110111000001010",
						 "000101110110110100111010",
						 "000101110110110001101010",
						 "000101110110101110011010",
						 "000101110110101011001010",
						 "000101110110100111111010",
						 "000101110110100100101010",
						 "000101110110100001011010",
						 "000101110110011110001010",
						 "000101110110011010111010",
						 "000101110110010111101010",
						 "000101110110010100011010",
						 "000101110111000101001010",
						 "000101110111000001111010",
						 "000101110110111110101010",
						 "000101110110111011011010",
						 "000101110110111000001010",
						 "000101110110110100111010",
						 "000101110110110001101010",
						 "000101110110101110011010",
						 "000101110110101011001010",
						 "000101110110100111111010",
						 "000101110110100100101010",
						 "000101110110100001011010",
						 "000101110110011110001010",
						 "000101110110011010111010",
						 "000101110110010111101010",
						 "000101110110010100011010",
						 "000101110111000101011001",
						 "000101110111000010001000",
						 "000101110110111110110111",
						 "000101110110111011100110",
						 "000101110110111000010101",
						 "000101110110110101000100",
						 "000101110110110001110011",
						 "000101110110101110100010",
						 "000101110110101011010001",
						 "000101110110101000000000",
						 "000101110110100100101111",
						 "000101110110100001011110",
						 "000101110110011110001101",
						 "000101110110011010111100",
						 "000101110110010111101011",
						 "000101110110010100011010",
						 "000101110100100010011011",
						 "000101110100011111001010",
						 "000101110100011011111001",
						 "000101110100011000101000",
						 "000101110100010101010111",
						 "000101110100010010000110",
						 "000101110100001110110101",
						 "000101110100001011100100",
						 "000101110100001000010011",
						 "000101110100000101000010",
						 "000101110100000001110001",
						 "000101110011111110100000",
						 "000101110011111011001111",
						 "000101110011110111111110",
						 "000101110011110100101101",
						 "000101110011110001011100",
						 "000101110100100010011011",
						 "000101110100011111001010",
						 "000101110100011011111001",
						 "000101110100011000101000",
						 "000101110100010101010111",
						 "000101110100010010000110",
						 "000101110100001110110101",
						 "000101110100001011100100",
						 "000101110100001000010011",
						 "000101110100000101000010",
						 "000101110100000001110001",
						 "000101110011111110100000",
						 "000101110011111011001111",
						 "000101110011110111111110",
						 "000101110011110100101101",
						 "000101110011110001011100",
						 "000101110100100010011011",
						 "000101110100011111001010",
						 "000101110100011011111001",
						 "000101110100011000101000",
						 "000101110100010101010111",
						 "000101110100010010000110",
						 "000101110100001110110101",
						 "000101110100001011100100",
						 "000101110100001000010011",
						 "000101110100000101000010",
						 "000101110100000001110001",
						 "000101110011111110100000",
						 "000101110011111011001111",
						 "000101110011110111111110",
						 "000101110011110100101101",
						 "000101110011110001011100",
						 "000101110001111111011101",
						 "000101110001111100001100",
						 "000101110001111000111011",
						 "000101110001110101101010",
						 "000101110001110010011001",
						 "000101110001101111001000",
						 "000101110001101011110111",
						 "000101110001101000100110",
						 "000101110001100101010101",
						 "000101110001100010000100",
						 "000101110001011110110011",
						 "000101110001011011100010",
						 "000101110001011000010001",
						 "000101110001010101000000",
						 "000101110001010001101111",
						 "000101110001001110011110",
						 "000101110001111111101100",
						 "000101110001111100011010",
						 "000101110001111001001000",
						 "000101110001110101110110",
						 "000101110001110010100100",
						 "000101110001101111010010",
						 "000101110001101100000000",
						 "000101110001101000101110",
						 "000101110001100101011100",
						 "000101110001100010001010",
						 "000101110001011110111000",
						 "000101110001011011100110",
						 "000101110001011000010100",
						 "000101110001010101000010",
						 "000101110001010001110000",
						 "000101110001001110011110",
						 "000101110001111111101100",
						 "000101110001111100011010",
						 "000101110001111001001000",
						 "000101110001110101110110",
						 "000101110001110010100100",
						 "000101110001101111010010",
						 "000101110001101100000000",
						 "000101110001101000101110",
						 "000101110001100101011100",
						 "000101110001100010001010",
						 "000101110001011110111000",
						 "000101110001011011100110",
						 "000101110001011000010100",
						 "000101110001010101000010",
						 "000101110001010001110000",
						 "000101110001001110011110",
						 "000101101111011100101110",
						 "000101101111011001011100",
						 "000101101111010110001010",
						 "000101101111010010111000",
						 "000101101111001111100110",
						 "000101101111001100010100",
						 "000101101111001001000010",
						 "000101101111000101110000",
						 "000101101111000010011110",
						 "000101101110111111001100",
						 "000101101110111011111010",
						 "000101101110111000101000",
						 "000101101110110101010110",
						 "000101101110110010000100",
						 "000101101110101110110010",
						 "000101101110101011100000",
						 "000101101111011100101110",
						 "000101101111011001011100",
						 "000101101111010110001010",
						 "000101101111010010111000",
						 "000101101111001111100110",
						 "000101101111001100010100",
						 "000101101111001001000010",
						 "000101101111000101110000",
						 "000101101111000010011110",
						 "000101101110111111001100",
						 "000101101110111011111010",
						 "000101101110111000101000",
						 "000101101110110101010110",
						 "000101101110110010000100",
						 "000101101110101110110010",
						 "000101101110101011100000",
						 "000101101111011100111101",
						 "000101101111011001101010",
						 "000101101111010110010111",
						 "000101101111010011000100",
						 "000101101111001111110001",
						 "000101101111001100011110",
						 "000101101111001001001011",
						 "000101101111000101111000",
						 "000101101111000010100101",
						 "000101101110111111010010",
						 "000101101110111011111111",
						 "000101101110111000101100",
						 "000101101110110101011001",
						 "000101101110110010000110",
						 "000101101110101110110011",
						 "000101101110101011100000",
						 "000101101100111001111111",
						 "000101101100110110101100",
						 "000101101100110011011001",
						 "000101101100110000000110",
						 "000101101100101100110011",
						 "000101101100101001100000",
						 "000101101100100110001101",
						 "000101101100100010111010",
						 "000101101100011111100111",
						 "000101101100011100010100",
						 "000101101100011001000001",
						 "000101101100010101101110",
						 "000101101100010010011011",
						 "000101101100001111001000",
						 "000101101100001011110101",
						 "000101101100001000100010",
						 "000101101100111001111111",
						 "000101101100110110101100",
						 "000101101100110011011001",
						 "000101101100110000000110",
						 "000101101100101100110011",
						 "000101101100101001100000",
						 "000101101100100110001101",
						 "000101101100100010111010",
						 "000101101100011111100111",
						 "000101101100011100010100",
						 "000101101100011001000001",
						 "000101101100010101101110",
						 "000101101100010010011011",
						 "000101101100001111001000",
						 "000101101100001011110101",
						 "000101101100001000100010",
						 "000101101100111001111111",
						 "000101101100110110101100",
						 "000101101100110011011001",
						 "000101101100110000000110",
						 "000101101100101100110011",
						 "000101101100101001100000",
						 "000101101100100110001101",
						 "000101101100100010111010",
						 "000101101100011111100111",
						 "000101101100011100010100",
						 "000101101100011001000001",
						 "000101101100010101101110",
						 "000101101100010010011011",
						 "000101101100001111001000",
						 "000101101100001011110101",
						 "000101101100001000100010",
						 "000101101010010111000001",
						 "000101101010010011101110",
						 "000101101010010000011011",
						 "000101101010001101001000",
						 "000101101010001001110101",
						 "000101101010000110100010",
						 "000101101010000011001111",
						 "000101101001111111111100",
						 "000101101001111100101001",
						 "000101101001111001010110",
						 "000101101001110110000011",
						 "000101101001110010110000",
						 "000101101001101111011101",
						 "000101101001101100001010",
						 "000101101001101000110111",
						 "000101101001100101100100",
						 "000101101010010111010000",
						 "000101101010010011111100",
						 "000101101010010000101000",
						 "000101101010001101010100",
						 "000101101010001010000000",
						 "000101101010000110101100",
						 "000101101010000011011000",
						 "000101101010000000000100",
						 "000101101001111100110000",
						 "000101101001111001011100",
						 "000101101001110110001000",
						 "000101101001110010110100",
						 "000101101001101111100000",
						 "000101101001101100001100",
						 "000101101001101000111000",
						 "000101101001100101100100",
						 "000101101010010111010000",
						 "000101101010010011111100",
						 "000101101010010000101000",
						 "000101101010001101010100",
						 "000101101010001010000000",
						 "000101101010000110101100",
						 "000101101010000011011000",
						 "000101101010000000000100",
						 "000101101001111100110000",
						 "000101101001111001011100",
						 "000101101001110110001000",
						 "000101101001110010110100",
						 "000101101001101111100000",
						 "000101101001101100001100",
						 "000101101001101000111000",
						 "000101101001100101100100",
						 "000101100111110100010010",
						 "000101100111110000111110",
						 "000101100111101101101010",
						 "000101100111101010010110",
						 "000101100111100111000010",
						 "000101100111100011101110",
						 "000101100111100000011010",
						 "000101100111011101000110",
						 "000101100111011001110010",
						 "000101100111010110011110",
						 "000101100111010011001010",
						 "000101100111001111110110",
						 "000101100111001100100010",
						 "000101100111001001001110",
						 "000101100111000101111010",
						 "000101100111000010100110",
						 "000101100111110100010010",
						 "000101100111110000111110",
						 "000101100111101101101010",
						 "000101100111101010010110",
						 "000101100111100111000010",
						 "000101100111100011101110",
						 "000101100111100000011010",
						 "000101100111011101000110",
						 "000101100111011001110010",
						 "000101100111010110011110",
						 "000101100111010011001010",
						 "000101100111001111110110",
						 "000101100111001100100010",
						 "000101100111001001001110",
						 "000101100111000101111010",
						 "000101100111000010100110",
						 "000101100111110100100001",
						 "000101100111110001001100",
						 "000101100111101101110111",
						 "000101100111101010100010",
						 "000101100111100111001101",
						 "000101100111100011111000",
						 "000101100111100000100011",
						 "000101100111011101001110",
						 "000101100111011001111001",
						 "000101100111010110100100",
						 "000101100111010011001111",
						 "000101100111001111111010",
						 "000101100111001100100101",
						 "000101100111001001010000",
						 "000101100111000101111011",
						 "000101100111000010100110",
						 "000101100101010001100011",
						 "000101100101001110001110",
						 "000101100101001010111001",
						 "000101100101000111100100",
						 "000101100101000100001111",
						 "000101100101000000111010",
						 "000101100100111101100101",
						 "000101100100111010010000",
						 "000101100100110110111011",
						 "000101100100110011100110",
						 "000101100100110000010001",
						 "000101100100101100111100",
						 "000101100100101001100111",
						 "000101100100100110010010",
						 "000101100100100010111101",
						 "000101100100011111101000",
						 "000101100101010001100011",
						 "000101100101001110001110",
						 "000101100101001010111001",
						 "000101100101000111100100",
						 "000101100101000100001111",
						 "000101100101000000111010",
						 "000101100100111101100101",
						 "000101100100111010010000",
						 "000101100100110110111011",
						 "000101100100110011100110",
						 "000101100100110000010001",
						 "000101100100101100111100",
						 "000101100100101001100111",
						 "000101100100100110010010",
						 "000101100100100010111101",
						 "000101100100011111101000",
						 "000101100101010001100011",
						 "000101100101001110001110",
						 "000101100101001010111001",
						 "000101100101000111100100",
						 "000101100101000100001111",
						 "000101100101000000111010",
						 "000101100100111101100101",
						 "000101100100111010010000",
						 "000101100100110110111011",
						 "000101100100110011100110",
						 "000101100100110000010001",
						 "000101100100101100111100",
						 "000101100100101001100111",
						 "000101100100100110010010",
						 "000101100100100010111101",
						 "000101100100011111101000",
						 "000101100010101110100101",
						 "000101100010101011010000",
						 "000101100010100111111011",
						 "000101100010100100100110",
						 "000101100010100001010001",
						 "000101100010011101111100",
						 "000101100010011010100111",
						 "000101100010010111010010",
						 "000101100010010011111101",
						 "000101100010010000101000",
						 "000101100010001101010011",
						 "000101100010001001111110",
						 "000101100010000110101001",
						 "000101100010000011010100",
						 "000101100001111111111111",
						 "000101100001111100101010",
						 "000101100010101110110100",
						 "000101100010101011011110",
						 "000101100010101000001000",
						 "000101100010100100110010",
						 "000101100010100001011100",
						 "000101100010011110000110",
						 "000101100010011010110000",
						 "000101100010010111011010",
						 "000101100010010100000100",
						 "000101100010010000101110",
						 "000101100010001101011000",
						 "000101100010001010000010",
						 "000101100010000110101100",
						 "000101100010000011010110",
						 "000101100010000000000000",
						 "000101100001111100101010",
						 "000101100010101110110100",
						 "000101100010101011011110",
						 "000101100010101000001000",
						 "000101100010100100110010",
						 "000101100010100001011100",
						 "000101100010011110000110",
						 "000101100010011010110000",
						 "000101100010010111011010",
						 "000101100010010100000100",
						 "000101100010010000101110",
						 "000101100010001101011000",
						 "000101100010001010000010",
						 "000101100010000110101100",
						 "000101100010000011010110",
						 "000101100010000000000000",
						 "000101100001111100101010",
						 "000101100000001011110110",
						 "000101100000001000100000",
						 "000101100000000101001010",
						 "000101100000000001110100",
						 "000101011111111110011110",
						 "000101011111111011001000",
						 "000101011111110111110010",
						 "000101011111110100011100",
						 "000101011111110001000110",
						 "000101011111101101110000",
						 "000101011111101010011010",
						 "000101011111100111000100",
						 "000101011111100011101110",
						 "000101011111100000011000",
						 "000101011111011101000010",
						 "000101011111011001101100",
						 "000101100000001011110110",
						 "000101100000001000100000",
						 "000101100000000101001010",
						 "000101100000000001110100",
						 "000101011111111110011110",
						 "000101011111111011001000",
						 "000101011111110111110010",
						 "000101011111110100011100",
						 "000101011111110001000110",
						 "000101011111101101110000",
						 "000101011111101010011010",
						 "000101011111100111000100",
						 "000101011111100011101110",
						 "000101011111100000011000",
						 "000101011111011101000010",
						 "000101011111011001101100",
						 "000101100000001011110110",
						 "000101100000001000100000",
						 "000101100000000101001010",
						 "000101100000000001110100",
						 "000101011111111110011110",
						 "000101011111111011001000",
						 "000101011111110111110010",
						 "000101011111110100011100",
						 "000101011111110001000110",
						 "000101011111101101110000",
						 "000101011111101010011010",
						 "000101011111100111000100",
						 "000101011111100011101110",
						 "000101011111100000011000",
						 "000101011111011101000010",
						 "000101011111011001101100",
						 "000101011101101001000111",
						 "000101011101100101110000",
						 "000101011101100010011001",
						 "000101011101011111000010",
						 "000101011101011011101011",
						 "000101011101011000010100",
						 "000101011101010100111101",
						 "000101011101010001100110",
						 "000101011101001110001111",
						 "000101011101001010111000",
						 "000101011101000111100001",
						 "000101011101000100001010",
						 "000101011101000000110011",
						 "000101011100111101011100",
						 "000101011100111010000101",
						 "000101011100110110101110",
						 "000101011101101001000111",
						 "000101011101100101110000",
						 "000101011101100010011001",
						 "000101011101011111000010",
						 "000101011101011011101011",
						 "000101011101011000010100",
						 "000101011101010100111101",
						 "000101011101010001100110",
						 "000101011101001110001111",
						 "000101011101001010111000",
						 "000101011101000111100001",
						 "000101011101000100001010",
						 "000101011101000000110011",
						 "000101011100111101011100",
						 "000101011100111010000101",
						 "000101011100110110101110",
						 "000101011101101001000111",
						 "000101011101100101110000",
						 "000101011101100010011001",
						 "000101011101011111000010",
						 "000101011101011011101011",
						 "000101011101011000010100",
						 "000101011101010100111101",
						 "000101011101010001100110",
						 "000101011101001110001111",
						 "000101011101001010111000",
						 "000101011101000111100001",
						 "000101011101000100001010",
						 "000101011101000000110011",
						 "000101011100111101011100",
						 "000101011100111010000101",
						 "000101011100110110101110",
						 "000101011011000110001001",
						 "000101011011000010110010",
						 "000101011010111111011011",
						 "000101011010111100000100",
						 "000101011010111000101101",
						 "000101011010110101010110",
						 "000101011010110001111111",
						 "000101011010101110101000",
						 "000101011010101011010001",
						 "000101011010100111111010",
						 "000101011010100100100011",
						 "000101011010100001001100",
						 "000101011010011101110101",
						 "000101011010011010011110",
						 "000101011010010111000111",
						 "000101011010010011110000",
						 "000101011011000110011000",
						 "000101011011000011000000",
						 "000101011010111111101000",
						 "000101011010111100010000",
						 "000101011010111000111000",
						 "000101011010110101100000",
						 "000101011010110010001000",
						 "000101011010101110110000",
						 "000101011010101011011000",
						 "000101011010101000000000",
						 "000101011010100100101000",
						 "000101011010100001010000",
						 "000101011010011101111000",
						 "000101011010011010100000",
						 "000101011010010111001000",
						 "000101011010010011110000",
						 "000101011011000110011000",
						 "000101011011000011000000",
						 "000101011010111111101000",
						 "000101011010111100010000",
						 "000101011010111000111000",
						 "000101011010110101100000",
						 "000101011010110010001000",
						 "000101011010101110110000",
						 "000101011010101011011000",
						 "000101011010101000000000",
						 "000101011010100100101000",
						 "000101011010100001010000",
						 "000101011010011101111000",
						 "000101011010011010100000",
						 "000101011010010111001000",
						 "000101011010010011110000",
						 "000101011000100011011010",
						 "000101011000100000000010",
						 "000101011000011100101010",
						 "000101011000011001010010",
						 "000101011000010101111010",
						 "000101011000010010100010",
						 "000101011000001111001010",
						 "000101011000001011110010",
						 "000101011000001000011010",
						 "000101011000000101000010",
						 "000101011000000001101010",
						 "000101010111111110010010",
						 "000101010111111010111010",
						 "000101010111110111100010",
						 "000101010111110100001010",
						 "000101010111110000110010",
						 "000101011000100011011010",
						 "000101011000100000000010",
						 "000101011000011100101010",
						 "000101011000011001010010",
						 "000101011000010101111010",
						 "000101011000010010100010",
						 "000101011000001111001010",
						 "000101011000001011110010",
						 "000101011000001000011010",
						 "000101011000000101000010",
						 "000101011000000001101010",
						 "000101010111111110010010",
						 "000101010111111010111010",
						 "000101010111110111100010",
						 "000101010111110100001010",
						 "000101010111110000110010",
						 "000101011000100011011010",
						 "000101011000100000000010",
						 "000101011000011100101010",
						 "000101011000011001010010",
						 "000101011000010101111010",
						 "000101011000010010100010",
						 "000101011000001111001010",
						 "000101011000001011110010",
						 "000101011000001000011010",
						 "000101011000000101000010",
						 "000101011000000001101010",
						 "000101010111111110010010",
						 "000101010111111010111010",
						 "000101010111110111100010",
						 "000101010111110100001010",
						 "000101010111110000110010",
						 "000101010110000000101011",
						 "000101010101111101010010",
						 "000101010101111001111001",
						 "000101010101110110100000",
						 "000101010101110011000111",
						 "000101010101101111101110",
						 "000101010101101100010101",
						 "000101010101101000111100",
						 "000101010101100101100011",
						 "000101010101100010001010",
						 "000101010101011110110001",
						 "000101010101011011011000",
						 "000101010101010111111111",
						 "000101010101010100100110",
						 "000101010101010001001101",
						 "000101010101001101110100",
						 "000101010110000000101011",
						 "000101010101111101010010",
						 "000101010101111001111001",
						 "000101010101110110100000",
						 "000101010101110011000111",
						 "000101010101101111101110",
						 "000101010101101100010101",
						 "000101010101101000111100",
						 "000101010101100101100011",
						 "000101010101100010001010",
						 "000101010101011110110001",
						 "000101010101011011011000",
						 "000101010101010111111111",
						 "000101010101010100100110",
						 "000101010101010001001101",
						 "000101010101001101110100",
						 "000101010110000000101011",
						 "000101010101111101010010",
						 "000101010101111001111001",
						 "000101010101110110100000",
						 "000101010101110011000111",
						 "000101010101101111101110",
						 "000101010101101100010101",
						 "000101010101101000111100",
						 "000101010101100101100011",
						 "000101010101100010001010",
						 "000101010101011110110001",
						 "000101010101011011011000",
						 "000101010101010111111111",
						 "000101010101010100100110",
						 "000101010101010001001101",
						 "000101010101001101110100",
						 "000101010011011101101101",
						 "000101010011011010010100",
						 "000101010011010110111011",
						 "000101010011010011100010",
						 "000101010011010000001001",
						 "000101010011001100110000",
						 "000101010011001001010111",
						 "000101010011000101111110",
						 "000101010011000010100101",
						 "000101010010111111001100",
						 "000101010010111011110011",
						 "000101010010111000011010",
						 "000101010010110101000001",
						 "000101010010110001101000",
						 "000101010010101110001111",
						 "000101010010101010110110",
						 "000101010011011101101101",
						 "000101010011011010010100",
						 "000101010011010110111011",
						 "000101010011010011100010",
						 "000101010011010000001001",
						 "000101010011001100110000",
						 "000101010011001001010111",
						 "000101010011000101111110",
						 "000101010011000010100101",
						 "000101010010111111001100",
						 "000101010010111011110011",
						 "000101010010111000011010",
						 "000101010010110101000001",
						 "000101010010110001101000",
						 "000101010010101110001111",
						 "000101010010101010110110",
						 "000101010011011101111100",
						 "000101010011011010100010",
						 "000101010011010111001000",
						 "000101010011010011101110",
						 "000101010011010000010100",
						 "000101010011001100111010",
						 "000101010011001001100000",
						 "000101010011000110000110",
						 "000101010011000010101100",
						 "000101010010111111010010",
						 "000101010010111011111000",
						 "000101010010111000011110",
						 "000101010010110101000100",
						 "000101010010110001101010",
						 "000101010010101110010000",
						 "000101010010101010110110",
						 "000101010000111010111110",
						 "000101010000110111100100",
						 "000101010000110100001010",
						 "000101010000110000110000",
						 "000101010000101101010110",
						 "000101010000101001111100",
						 "000101010000100110100010",
						 "000101010000100011001000",
						 "000101010000011111101110",
						 "000101010000011100010100",
						 "000101010000011000111010",
						 "000101010000010101100000",
						 "000101010000010010000110",
						 "000101010000001110101100",
						 "000101010000001011010010",
						 "000101010000000111111000",
						 "000101010000111010111110",
						 "000101010000110111100100",
						 "000101010000110100001010",
						 "000101010000110000110000",
						 "000101010000101101010110",
						 "000101010000101001111100",
						 "000101010000100110100010",
						 "000101010000100011001000",
						 "000101010000011111101110",
						 "000101010000011100010100",
						 "000101010000011000111010",
						 "000101010000010101100000",
						 "000101010000010010000110",
						 "000101010000001110101100",
						 "000101010000001011010010",
						 "000101010000000111111000",
						 "000101010000111010111110",
						 "000101010000110111100100",
						 "000101010000110100001010",
						 "000101010000110000110000",
						 "000101010000101101010110",
						 "000101010000101001111100",
						 "000101010000100110100010",
						 "000101010000100011001000",
						 "000101010000011111101110",
						 "000101010000011100010100",
						 "000101010000011000111010",
						 "000101010000010101100000",
						 "000101010000010010000110",
						 "000101010000001110101100",
						 "000101010000001011010010",
						 "000101010000000111111000",
						 "000101001110011000000000",
						 "000101001110010100100110",
						 "000101001110010001001100",
						 "000101001110001101110010",
						 "000101001110001010011000",
						 "000101001110000110111110",
						 "000101001110000011100100",
						 "000101001110000000001010",
						 "000101001101111100110000",
						 "000101001101111001010110",
						 "000101001101110101111100",
						 "000101001101110010100010",
						 "000101001101101111001000",
						 "000101001101101011101110",
						 "000101001101101000010100",
						 "000101001101100100111010",
						 "000101001110011000001111",
						 "000101001110010100110100",
						 "000101001110010001011001",
						 "000101001110001101111110",
						 "000101001110001010100011",
						 "000101001110000111001000",
						 "000101001110000011101101",
						 "000101001110000000010010",
						 "000101001101111100110111",
						 "000101001101111001011100",
						 "000101001101110110000001",
						 "000101001101110010100110",
						 "000101001101101111001011",
						 "000101001101101011110000",
						 "000101001101101000010101",
						 "000101001101100100111010",
						 "000101001110011000001111",
						 "000101001110010100110100",
						 "000101001110010001011001",
						 "000101001110001101111110",
						 "000101001110001010100011",
						 "000101001110000111001000",
						 "000101001110000011101101",
						 "000101001110000000010010",
						 "000101001101111100110111",
						 "000101001101111001011100",
						 "000101001101110110000001",
						 "000101001101110010100110",
						 "000101001101101111001011",
						 "000101001101101011110000",
						 "000101001101101000010101",
						 "000101001101100100111010",
						 "000101001011110101010001",
						 "000101001011110001110110",
						 "000101001011101110011011",
						 "000101001011101011000000",
						 "000101001011100111100101",
						 "000101001011100100001010",
						 "000101001011100000101111",
						 "000101001011011101010100",
						 "000101001011011001111001",
						 "000101001011010110011110",
						 "000101001011010011000011",
						 "000101001011001111101000",
						 "000101001011001100001101",
						 "000101001011001000110010",
						 "000101001011000101010111",
						 "000101001011000001111100",
						 "000101001011110101010001",
						 "000101001011110001110110",
						 "000101001011101110011011",
						 "000101001011101011000000",
						 "000101001011100111100101",
						 "000101001011100100001010",
						 "000101001011100000101111",
						 "000101001011011101010100",
						 "000101001011011001111001",
						 "000101001011010110011110",
						 "000101001011010011000011",
						 "000101001011001111101000",
						 "000101001011001100001101",
						 "000101001011001000110010",
						 "000101001011000101010111",
						 "000101001011000001111100",
						 "000101001011110101010001",
						 "000101001011110001110110",
						 "000101001011101110011011",
						 "000101001011101011000000",
						 "000101001011100111100101",
						 "000101001011100100001010",
						 "000101001011100000101111",
						 "000101001011011101010100",
						 "000101001011011001111001",
						 "000101001011010110011110",
						 "000101001011010011000011",
						 "000101001011001111101000",
						 "000101001011001100001101",
						 "000101001011001000110010",
						 "000101001011000101010111",
						 "000101001011000001111100",
						 "000101001001010010100010",
						 "000101001001001111000110",
						 "000101001001001011101010",
						 "000101001001001000001110",
						 "000101001001000100110010",
						 "000101001001000001010110",
						 "000101001000111101111010",
						 "000101001000111010011110",
						 "000101001000110111000010",
						 "000101001000110011100110",
						 "000101001000110000001010",
						 "000101001000101100101110",
						 "000101001000101001010010",
						 "000101001000100101110110",
						 "000101001000100010011010",
						 "000101001000011110111110",
						 "000101001001010010100010",
						 "000101001001001111000110",
						 "000101001001001011101010",
						 "000101001001001000001110",
						 "000101001001000100110010",
						 "000101001001000001010110",
						 "000101001000111101111010",
						 "000101001000111010011110",
						 "000101001000110111000010",
						 "000101001000110011100110",
						 "000101001000110000001010",
						 "000101001000101100101110",
						 "000101001000101001010010",
						 "000101001000100101110110",
						 "000101001000100010011010",
						 "000101001000011110111110",
						 "000101001001010010100010",
						 "000101001001001111000110",
						 "000101001001001011101010",
						 "000101001001001000001110",
						 "000101001001000100110010",
						 "000101001001000001010110",
						 "000101001000111101111010",
						 "000101001000111010011110",
						 "000101001000110111000010",
						 "000101001000110011100110",
						 "000101001000110000001010",
						 "000101001000101100101110",
						 "000101001000101001010010",
						 "000101001000100101110110",
						 "000101001000100010011010",
						 "000101001000011110111110",
						 "000101000110101111100100",
						 "000101000110101100001000",
						 "000101000110101000101100",
						 "000101000110100101010000",
						 "000101000110100001110100",
						 "000101000110011110011000",
						 "000101000110011010111100",
						 "000101000110010111100000",
						 "000101000110010100000100",
						 "000101000110010000101000",
						 "000101000110001101001100",
						 "000101000110001001110000",
						 "000101000110000110010100",
						 "000101000110000010111000",
						 "000101000101111111011100",
						 "000101000101111100000000",
						 "000101000110101111100100",
						 "000101000110101100001000",
						 "000101000110101000101100",
						 "000101000110100101010000",
						 "000101000110100001110100",
						 "000101000110011110011000",
						 "000101000110011010111100",
						 "000101000110010111100000",
						 "000101000110010100000100",
						 "000101000110010000101000",
						 "000101000110001101001100",
						 "000101000110001001110000",
						 "000101000110000110010100",
						 "000101000110000010111000",
						 "000101000101111111011100",
						 "000101000101111100000000",
						 "000101000110101111110011",
						 "000101000110101100010110",
						 "000101000110101000111001",
						 "000101000110100101011100",
						 "000101000110100001111111",
						 "000101000110011110100010",
						 "000101000110011011000101",
						 "000101000110010111101000",
						 "000101000110010100001011",
						 "000101000110010000101110",
						 "000101000110001101010001",
						 "000101000110001001110100",
						 "000101000110000110010111",
						 "000101000110000010111010",
						 "000101000101111111011101",
						 "000101000101111100000000",
						 "000101000100001100110101",
						 "000101000100001001011000",
						 "000101000100000101111011",
						 "000101000100000010011110",
						 "000101000011111111000001",
						 "000101000011111011100100",
						 "000101000011111000000111",
						 "000101000011110100101010",
						 "000101000011110001001101",
						 "000101000011101101110000",
						 "000101000011101010010011",
						 "000101000011100110110110",
						 "000101000011100011011001",
						 "000101000011011111111100",
						 "000101000011011100011111",
						 "000101000011011001000010",
						 "000101000100001100110101",
						 "000101000100001001011000",
						 "000101000100000101111011",
						 "000101000100000010011110",
						 "000101000011111111000001",
						 "000101000011111011100100",
						 "000101000011111000000111",
						 "000101000011110100101010",
						 "000101000011110001001101",
						 "000101000011101101110000",
						 "000101000011101010010011",
						 "000101000011100110110110",
						 "000101000011100011011001",
						 "000101000011011111111100",
						 "000101000011011100011111",
						 "000101000011011001000010",
						 "000101000100001100110101",
						 "000101000100001001011000",
						 "000101000100000101111011",
						 "000101000100000010011110",
						 "000101000011111111000001",
						 "000101000011111011100100",
						 "000101000011111000000111",
						 "000101000011110100101010",
						 "000101000011110001001101",
						 "000101000011101101110000",
						 "000101000011101010010011",
						 "000101000011100110110110",
						 "000101000011100011011001",
						 "000101000011011111111100",
						 "000101000011011100011111",
						 "000101000011011001000010",
						 "000101000001101001110111",
						 "000101000001100110011010",
						 "000101000001100010111101",
						 "000101000001011111100000",
						 "000101000001011100000011",
						 "000101000001011000100110",
						 "000101000001010101001001",
						 "000101000001010001101100",
						 "000101000001001110001111",
						 "000101000001001010110010",
						 "000101000001000111010101",
						 "000101000001000011111000",
						 "000101000001000000011011",
						 "000101000000111100111110",
						 "000101000000111001100001",
						 "000101000000110110000100",
						 "000101000001101010000110",
						 "000101000001100110101000",
						 "000101000001100011001010",
						 "000101000001011111101100",
						 "000101000001011100001110",
						 "000101000001011000110000",
						 "000101000001010101010010",
						 "000101000001010001110100",
						 "000101000001001110010110",
						 "000101000001001010111000",
						 "000101000001000111011010",
						 "000101000001000011111100",
						 "000101000001000000011110",
						 "000101000000111101000000",
						 "000101000000111001100010",
						 "000101000000110110000100",
						 "000101000001101010000110",
						 "000101000001100110101000",
						 "000101000001100011001010",
						 "000101000001011111101100",
						 "000101000001011100001110",
						 "000101000001011000110000",
						 "000101000001010101010010",
						 "000101000001010001110100",
						 "000101000001001110010110",
						 "000101000001001010111000",
						 "000101000001000111011010",
						 "000101000001000011111100",
						 "000101000001000000011110",
						 "000101000000111101000000",
						 "000101000000111001100010",
						 "000101000000110110000100",
						 "000100111111000111001000",
						 "000100111111000011101010",
						 "000100111111000000001100",
						 "000100111110111100101110",
						 "000100111110111001010000",
						 "000100111110110101110010",
						 "000100111110110010010100",
						 "000100111110101110110110",
						 "000100111110101011011000",
						 "000100111110100111111010",
						 "000100111110100100011100",
						 "000100111110100000111110",
						 "000100111110011101100000",
						 "000100111110011010000010",
						 "000100111110010110100100",
						 "000100111110010011000110",
						 "000100111111000111001000",
						 "000100111111000011101010",
						 "000100111111000000001100",
						 "000100111110111100101110",
						 "000100111110111001010000",
						 "000100111110110101110010",
						 "000100111110110010010100",
						 "000100111110101110110110",
						 "000100111110101011011000",
						 "000100111110100111111010",
						 "000100111110100100011100",
						 "000100111110100000111110",
						 "000100111110011101100000",
						 "000100111110011010000010",
						 "000100111110010110100100",
						 "000100111110010011000110",
						 "000100111111000111001000",
						 "000100111111000011101010",
						 "000100111111000000001100",
						 "000100111110111100101110",
						 "000100111110111001010000",
						 "000100111110110101110010",
						 "000100111110110010010100",
						 "000100111110101110110110",
						 "000100111110101011011000",
						 "000100111110100111111010",
						 "000100111110100100011100",
						 "000100111110100000111110",
						 "000100111110011101100000",
						 "000100111110011010000010",
						 "000100111110010110100100",
						 "000100111110010011000110",
						 "000100111100100100011001",
						 "000100111100100000111010",
						 "000100111100011101011011",
						 "000100111100011001111100",
						 "000100111100010110011101",
						 "000100111100010010111110",
						 "000100111100001111011111",
						 "000100111100001100000000",
						 "000100111100001000100001",
						 "000100111100000101000010",
						 "000100111100000001100011",
						 "000100111011111110000100",
						 "000100111011111010100101",
						 "000100111011110111000110",
						 "000100111011110011100111",
						 "000100111011110000001000",
						 "000100111100100100011001",
						 "000100111100100000111010",
						 "000100111100011101011011",
						 "000100111100011001111100",
						 "000100111100010110011101",
						 "000100111100010010111110",
						 "000100111100001111011111",
						 "000100111100001100000000",
						 "000100111100001000100001",
						 "000100111100000101000010",
						 "000100111100000001100011",
						 "000100111011111110000100",
						 "000100111011111010100101",
						 "000100111011110111000110",
						 "000100111011110011100111",
						 "000100111011110000001000",
						 "000100111100100100011001",
						 "000100111100100000111010",
						 "000100111100011101011011",
						 "000100111100011001111100",
						 "000100111100010110011101",
						 "000100111100010010111110",
						 "000100111100001111011111",
						 "000100111100001100000000",
						 "000100111100001000100001",
						 "000100111100000101000010",
						 "000100111100000001100011",
						 "000100111011111110000100",
						 "000100111011111010100101",
						 "000100111011110111000110",
						 "000100111011110011100111",
						 "000100111011110000001000",
						 "000100111010000001011011",
						 "000100111001111101111100",
						 "000100111001111010011101",
						 "000100111001110110111110",
						 "000100111001110011011111",
						 "000100111001110000000000",
						 "000100111001101100100001",
						 "000100111001101001000010",
						 "000100111001100101100011",
						 "000100111001100010000100",
						 "000100111001011110100101",
						 "000100111001011011000110",
						 "000100111001010111100111",
						 "000100111001010100001000",
						 "000100111001010000101001",
						 "000100111001001101001010",
						 "000100111010000001011011",
						 "000100111001111101111100",
						 "000100111001111010011101",
						 "000100111001110110111110",
						 "000100111001110011011111",
						 "000100111001110000000000",
						 "000100111001101100100001",
						 "000100111001101001000010",
						 "000100111001100101100011",
						 "000100111001100010000100",
						 "000100111001011110100101",
						 "000100111001011011000110",
						 "000100111001010111100111",
						 "000100111001010100001000",
						 "000100111001010000101001",
						 "000100111001001101001010",
						 "000100111010000001011011",
						 "000100111001111101111100",
						 "000100111001111010011101",
						 "000100111001110110111110",
						 "000100111001110011011111",
						 "000100111001110000000000",
						 "000100111001101100100001",
						 "000100111001101001000010",
						 "000100111001100101100011",
						 "000100111001100010000100",
						 "000100111001011110100101",
						 "000100111001011011000110",
						 "000100111001010111100111",
						 "000100111001010100001000",
						 "000100111001010000101001",
						 "000100111001001101001010",
						 "000100110111011110101100",
						 "000100110111011011001100",
						 "000100110111010111101100",
						 "000100110111010100001100",
						 "000100110111010000101100",
						 "000100110111001101001100",
						 "000100110111001001101100",
						 "000100110111000110001100",
						 "000100110111000010101100",
						 "000100110110111111001100",
						 "000100110110111011101100",
						 "000100110110111000001100",
						 "000100110110110100101100",
						 "000100110110110001001100",
						 "000100110110101101101100",
						 "000100110110101010001100",
						 "000100110111011110101100",
						 "000100110111011011001100",
						 "000100110111010111101100",
						 "000100110111010100001100",
						 "000100110111010000101100",
						 "000100110111001101001100",
						 "000100110111001001101100",
						 "000100110111000110001100",
						 "000100110111000010101100",
						 "000100110110111111001100",
						 "000100110110111011101100",
						 "000100110110111000001100",
						 "000100110110110100101100",
						 "000100110110110001001100",
						 "000100110110101101101100",
						 "000100110110101010001100",
						 "000100110111011110101100",
						 "000100110111011011001100",
						 "000100110111010111101100",
						 "000100110111010100001100",
						 "000100110111010000101100",
						 "000100110111001101001100",
						 "000100110111001001101100",
						 "000100110111000110001100",
						 "000100110111000010101100",
						 "000100110110111111001100",
						 "000100110110111011101100",
						 "000100110110111000001100",
						 "000100110110110100101100",
						 "000100110110110001001100",
						 "000100110110101101101100",
						 "000100110110101010001100",
						 "000100110100111011101110",
						 "000100110100111000001110",
						 "000100110100110100101110",
						 "000100110100110001001110",
						 "000100110100101101101110",
						 "000100110100101010001110",
						 "000100110100100110101110",
						 "000100110100100011001110",
						 "000100110100011111101110",
						 "000100110100011100001110",
						 "000100110100011000101110",
						 "000100110100010101001110",
						 "000100110100010001101110",
						 "000100110100001110001110",
						 "000100110100001010101110",
						 "000100110100000111001110",
						 "000100110100111011101110",
						 "000100110100111000001110",
						 "000100110100110100101110",
						 "000100110100110001001110",
						 "000100110100101101101110",
						 "000100110100101010001110",
						 "000100110100100110101110",
						 "000100110100100011001110",
						 "000100110100011111101110",
						 "000100110100011100001110",
						 "000100110100011000101110",
						 "000100110100010101001110",
						 "000100110100010001101110",
						 "000100110100001110001110",
						 "000100110100001010101110",
						 "000100110100000111001110",
						 "000100110100111011111101",
						 "000100110100111000011100",
						 "000100110100110100111011",
						 "000100110100110001011010",
						 "000100110100101101111001",
						 "000100110100101010011000",
						 "000100110100100110110111",
						 "000100110100100011010110",
						 "000100110100011111110101",
						 "000100110100011100010100",
						 "000100110100011000110011",
						 "000100110100010101010010",
						 "000100110100010001110001",
						 "000100110100001110010000",
						 "000100110100001010101111",
						 "000100110100000111001110",
						 "000100110010011000111111",
						 "000100110010010101011110",
						 "000100110010010001111101",
						 "000100110010001110011100",
						 "000100110010001010111011",
						 "000100110010000111011010",
						 "000100110010000011111001",
						 "000100110010000000011000",
						 "000100110001111100110111",
						 "000100110001111001010110",
						 "000100110001110101110101",
						 "000100110001110010010100",
						 "000100110001101110110011",
						 "000100110001101011010010",
						 "000100110001100111110001",
						 "000100110001100100010000",
						 "000100110010011000111111",
						 "000100110010010101011110",
						 "000100110010010001111101",
						 "000100110010001110011100",
						 "000100110010001010111011",
						 "000100110010000111011010",
						 "000100110010000011111001",
						 "000100110010000000011000",
						 "000100110001111100110111",
						 "000100110001111001010110",
						 "000100110001110101110101",
						 "000100110001110010010100",
						 "000100110001101110110011",
						 "000100110001101011010010",
						 "000100110001100111110001",
						 "000100110001100100010000",
						 "000100110010011000111111",
						 "000100110010010101011110",
						 "000100110010010001111101",
						 "000100110010001110011100",
						 "000100110010001010111011",
						 "000100110010000111011010",
						 "000100110010000011111001",
						 "000100110010000000011000",
						 "000100110001111100110111",
						 "000100110001111001010110",
						 "000100110001110101110101",
						 "000100110001110010010100",
						 "000100110001101110110011",
						 "000100110001101011010010",
						 "000100110001100111110001",
						 "000100110001100100010000",
						 "000100101111110110000001",
						 "000100101111110010100000",
						 "000100101111101110111111",
						 "000100101111101011011110",
						 "000100101111100111111101",
						 "000100101111100100011100",
						 "000100101111100000111011",
						 "000100101111011101011010",
						 "000100101111011001111001",
						 "000100101111010110011000",
						 "000100101111010010110111",
						 "000100101111001111010110",
						 "000100101111001011110101",
						 "000100101111001000010100",
						 "000100101111000100110011",
						 "000100101111000001010010",
						 "000100101111110110010000",
						 "000100101111110010101110",
						 "000100101111101111001100",
						 "000100101111101011101010",
						 "000100101111101000001000",
						 "000100101111100100100110",
						 "000100101111100001000100",
						 "000100101111011101100010",
						 "000100101111011010000000",
						 "000100101111010110011110",
						 "000100101111010010111100",
						 "000100101111001111011010",
						 "000100101111001011111000",
						 "000100101111001000010110",
						 "000100101111000100110100",
						 "000100101111000001010010",
						 "000100101101010011010010",
						 "000100101101001111110000",
						 "000100101101001100001110",
						 "000100101101001000101100",
						 "000100101101000101001010",
						 "000100101101000001101000",
						 "000100101100111110000110",
						 "000100101100111010100100",
						 "000100101100110111000010",
						 "000100101100110011100000",
						 "000100101100101111111110",
						 "000100101100101100011100",
						 "000100101100101000111010",
						 "000100101100100101011000",
						 "000100101100100001110110",
						 "000100101100011110010100",
						 "000100101101010011010010",
						 "000100101101001111110000",
						 "000100101101001100001110",
						 "000100101101001000101100",
						 "000100101101000101001010",
						 "000100101101000001101000",
						 "000100101100111110000110",
						 "000100101100111010100100",
						 "000100101100110111000010",
						 "000100101100110011100000",
						 "000100101100101111111110",
						 "000100101100101100011100",
						 "000100101100101000111010",
						 "000100101100100101011000",
						 "000100101100100001110110",
						 "000100101100011110010100",
						 "000100101101010011010010",
						 "000100101101001111110000",
						 "000100101101001100001110",
						 "000100101101001000101100",
						 "000100101101000101001010",
						 "000100101101000001101000",
						 "000100101100111110000110",
						 "000100101100111010100100",
						 "000100101100110111000010",
						 "000100101100110011100000",
						 "000100101100101111111110",
						 "000100101100101100011100",
						 "000100101100101000111010",
						 "000100101100100101011000",
						 "000100101100100001110110",
						 "000100101100011110010100",
						 "000100101010110000010100",
						 "000100101010101100110010",
						 "000100101010101001010000",
						 "000100101010100101101110",
						 "000100101010100010001100",
						 "000100101010011110101010",
						 "000100101010011011001000",
						 "000100101010010111100110",
						 "000100101010010100000100",
						 "000100101010010000100010",
						 "000100101010001101000000",
						 "000100101010001001011110",
						 "000100101010000101111100",
						 "000100101010000010011010",
						 "000100101001111110111000",
						 "000100101001111011010110",
						 "000100101010110000010100",
						 "000100101010101100110010",
						 "000100101010101001010000",
						 "000100101010100101101110",
						 "000100101010100010001100",
						 "000100101010011110101010",
						 "000100101010011011001000",
						 "000100101010010111100110",
						 "000100101010010100000100",
						 "000100101010010000100010",
						 "000100101010001101000000",
						 "000100101010001001011110",
						 "000100101010000101111100",
						 "000100101010000010011010",
						 "000100101001111110111000",
						 "000100101001111011010110",
						 "000100101010110000100011",
						 "000100101010101101000000",
						 "000100101010101001011101",
						 "000100101010100101111010",
						 "000100101010100010010111",
						 "000100101010011110110100",
						 "000100101010011011010001",
						 "000100101010010111101110",
						 "000100101010010100001011",
						 "000100101010010000101000",
						 "000100101010001101000101",
						 "000100101010001001100010",
						 "000100101010000101111111",
						 "000100101010000010011100",
						 "000100101001111110111001",
						 "000100101001111011010110",
						 "000100101000001101100101",
						 "000100101000001010000010",
						 "000100101000000110011111",
						 "000100101000000010111100",
						 "000100100111111111011001",
						 "000100100111111011110110",
						 "000100100111111000010011",
						 "000100100111110100110000",
						 "000100100111110001001101",
						 "000100100111101101101010",
						 "000100100111101010000111",
						 "000100100111100110100100",
						 "000100100111100011000001",
						 "000100100111011111011110",
						 "000100100111011011111011",
						 "000100100111011000011000",
						 "000100101000001101100101",
						 "000100101000001010000010",
						 "000100101000000110011111",
						 "000100101000000010111100",
						 "000100100111111111011001",
						 "000100100111111011110110",
						 "000100100111111000010011",
						 "000100100111110100110000",
						 "000100100111110001001101",
						 "000100100111101101101010",
						 "000100100111101010000111",
						 "000100100111100110100100",
						 "000100100111100011000001",
						 "000100100111011111011110",
						 "000100100111011011111011",
						 "000100100111011000011000",
						 "000100101000001101100101",
						 "000100101000001010000010",
						 "000100101000000110011111",
						 "000100101000000010111100",
						 "000100100111111111011001",
						 "000100100111111011110110",
						 "000100100111111000010011",
						 "000100100111110100110000",
						 "000100100111110001001101",
						 "000100100111101101101010",
						 "000100100111101010000111",
						 "000100100111100110100100",
						 "000100100111100011000001",
						 "000100100111011111011110",
						 "000100100111011011111011",
						 "000100100111011000011000",
						 "000100100101101010100111",
						 "000100100101100111000100",
						 "000100100101100011100001",
						 "000100100101011111111110",
						 "000100100101011100011011",
						 "000100100101011000111000",
						 "000100100101010101010101",
						 "000100100101010001110010",
						 "000100100101001110001111",
						 "000100100101001010101100",
						 "000100100101000111001001",
						 "000100100101000011100110",
						 "000100100101000000000011",
						 "000100100100111100100000",
						 "000100100100111000111101",
						 "000100100100110101011010",
						 "000100100101101010110110",
						 "000100100101100111010010",
						 "000100100101100011101110",
						 "000100100101100000001010",
						 "000100100101011100100110",
						 "000100100101011001000010",
						 "000100100101010101011110",
						 "000100100101010001111010",
						 "000100100101001110010110",
						 "000100100101001010110010",
						 "000100100101000111001110",
						 "000100100101000011101010",
						 "000100100101000000000110",
						 "000100100100111100100010",
						 "000100100100111000111110",
						 "000100100100110101011010",
						 "000100100101101010110110",
						 "000100100101100111010010",
						 "000100100101100011101110",
						 "000100100101100000001010",
						 "000100100101011100100110",
						 "000100100101011001000010",
						 "000100100101010101011110",
						 "000100100101010001111010",
						 "000100100101001110010110",
						 "000100100101001010110010",
						 "000100100101000111001110",
						 "000100100101000011101010",
						 "000100100101000000000110",
						 "000100100100111100100010",
						 "000100100100111000111110",
						 "000100100100110101011010",
						 "000100100011000111111000",
						 "000100100011000100010100",
						 "000100100011000000110000",
						 "000100100010111101001100",
						 "000100100010111001101000",
						 "000100100010110110000100",
						 "000100100010110010100000",
						 "000100100010101110111100",
						 "000100100010101011011000",
						 "000100100010100111110100",
						 "000100100010100100010000",
						 "000100100010100000101100",
						 "000100100010011101001000",
						 "000100100010011001100100",
						 "000100100010010110000000",
						 "000100100010010010011100",
						 "000100100011000111111000",
						 "000100100011000100010100",
						 "000100100011000000110000",
						 "000100100010111101001100",
						 "000100100010111001101000",
						 "000100100010110110000100",
						 "000100100010110010100000",
						 "000100100010101110111100",
						 "000100100010101011011000",
						 "000100100010100111110100",
						 "000100100010100100010000",
						 "000100100010100000101100",
						 "000100100010011101001000",
						 "000100100010011001100100",
						 "000100100010010110000000",
						 "000100100010010010011100",
						 "000100100011000111111000",
						 "000100100011000100010100",
						 "000100100011000000110000",
						 "000100100010111101001100",
						 "000100100010111001101000",
						 "000100100010110110000100",
						 "000100100010110010100000",
						 "000100100010101110111100",
						 "000100100010101011011000",
						 "000100100010100111110100",
						 "000100100010100100010000",
						 "000100100010100000101100",
						 "000100100010011101001000",
						 "000100100010011001100100",
						 "000100100010010110000000",
						 "000100100010010010011100",
						 "000100100000100100111010",
						 "000100100000100001010110",
						 "000100100000011101110010",
						 "000100100000011010001110",
						 "000100100000010110101010",
						 "000100100000010011000110",
						 "000100100000001111100010",
						 "000100100000001011111110",
						 "000100100000001000011010",
						 "000100100000000100110110",
						 "000100100000000001010010",
						 "000100011111111101101110",
						 "000100011111111010001010",
						 "000100011111110110100110",
						 "000100011111110011000010",
						 "000100011111101111011110",
						 "000100100000100101001001",
						 "000100100000100001100100",
						 "000100100000011101111111",
						 "000100100000011010011010",
						 "000100100000010110110101",
						 "000100100000010011010000",
						 "000100100000001111101011",
						 "000100100000001100000110",
						 "000100100000001000100001",
						 "000100100000000100111100",
						 "000100100000000001010111",
						 "000100011111111101110010",
						 "000100011111111010001101",
						 "000100011111110110101000",
						 "000100011111110011000011",
						 "000100011111101111011110",
						 "000100100000100101001001",
						 "000100100000100001100100",
						 "000100100000011101111111",
						 "000100100000011010011010",
						 "000100100000010110110101",
						 "000100100000010011010000",
						 "000100100000001111101011",
						 "000100100000001100000110",
						 "000100100000001000100001",
						 "000100100000000100111100",
						 "000100100000000001010111",
						 "000100011111111101110010",
						 "000100011111111010001101",
						 "000100011111110110101000",
						 "000100011111110011000011",
						 "000100011111101111011110",
						 "000100011110000010001011",
						 "000100011101111110100110",
						 "000100011101111011000001",
						 "000100011101110111011100",
						 "000100011101110011110111",
						 "000100011101110000010010",
						 "000100011101101100101101",
						 "000100011101101001001000",
						 "000100011101100101100011",
						 "000100011101100001111110",
						 "000100011101011110011001",
						 "000100011101011010110100",
						 "000100011101010111001111",
						 "000100011101010011101010",
						 "000100011101010000000101",
						 "000100011101001100100000",
						 "000100011110000010001011",
						 "000100011101111110100110",
						 "000100011101111011000001",
						 "000100011101110111011100",
						 "000100011101110011110111",
						 "000100011101110000010010",
						 "000100011101101100101101",
						 "000100011101101001001000",
						 "000100011101100101100011",
						 "000100011101100001111110",
						 "000100011101011110011001",
						 "000100011101011010110100",
						 "000100011101010111001111",
						 "000100011101010011101010",
						 "000100011101010000000101",
						 "000100011101001100100000",
						 "000100011011011111001101",
						 "000100011011011011101000",
						 "000100011011011000000011",
						 "000100011011010100011110",
						 "000100011011010000111001",
						 "000100011011001101010100",
						 "000100011011001001101111",
						 "000100011011000110001010",
						 "000100011011000010100101",
						 "000100011010111111000000",
						 "000100011010111011011011",
						 "000100011010110111110110",
						 "000100011010110100010001",
						 "000100011010110000101100",
						 "000100011010101101000111",
						 "000100011010101001100010",
						 "000100011011011111001101",
						 "000100011011011011101000",
						 "000100011011011000000011",
						 "000100011011010100011110",
						 "000100011011010000111001",
						 "000100011011001101010100",
						 "000100011011001001101111",
						 "000100011011000110001010",
						 "000100011011000010100101",
						 "000100011010111111000000",
						 "000100011010111011011011",
						 "000100011010110111110110",
						 "000100011010110100010001",
						 "000100011010110000101100",
						 "000100011010101101000111",
						 "000100011010101001100010",
						 "000100011011011111011100",
						 "000100011011011011110110",
						 "000100011011011000010000",
						 "000100011011010100101010",
						 "000100011011010001000100",
						 "000100011011001101011110",
						 "000100011011001001111000",
						 "000100011011000110010010",
						 "000100011011000010101100",
						 "000100011010111111000110",
						 "000100011010111011100000",
						 "000100011010110111111010",
						 "000100011010110100010100",
						 "000100011010110000101110",
						 "000100011010101101001000",
						 "000100011010101001100010",
						 "000100011000111100011110",
						 "000100011000111000111000",
						 "000100011000110101010010",
						 "000100011000110001101100",
						 "000100011000101110000110",
						 "000100011000101010100000",
						 "000100011000100110111010",
						 "000100011000100011010100",
						 "000100011000011111101110",
						 "000100011000011100001000",
						 "000100011000011000100010",
						 "000100011000010100111100",
						 "000100011000010001010110",
						 "000100011000001101110000",
						 "000100011000001010001010",
						 "000100011000000110100100",
						 "000100011000111100011110",
						 "000100011000111000111000",
						 "000100011000110101010010",
						 "000100011000110001101100",
						 "000100011000101110000110",
						 "000100011000101010100000",
						 "000100011000100110111010",
						 "000100011000100011010100",
						 "000100011000011111101110",
						 "000100011000011100001000",
						 "000100011000011000100010",
						 "000100011000010100111100",
						 "000100011000010001010110",
						 "000100011000001101110000",
						 "000100011000001010001010",
						 "000100011000000110100100",
						 "000100011000111100011110",
						 "000100011000111000111000",
						 "000100011000110101010010",
						 "000100011000110001101100",
						 "000100011000101110000110",
						 "000100011000101010100000",
						 "000100011000100110111010",
						 "000100011000100011010100",
						 "000100011000011111101110",
						 "000100011000011100001000",
						 "000100011000011000100010",
						 "000100011000010100111100",
						 "000100011000010001010110",
						 "000100011000001101110000",
						 "000100011000001010001010",
						 "000100011000000110100100",
						 "000100010110011001100000",
						 "000100010110010101111010",
						 "000100010110010010010100",
						 "000100010110001110101110",
						 "000100010110001011001000",
						 "000100010110000111100010",
						 "000100010110000011111100",
						 "000100010110000000010110",
						 "000100010101111100110000",
						 "000100010101111001001010",
						 "000100010101110101100100",
						 "000100010101110001111110",
						 "000100010101101110011000",
						 "000100010101101010110010",
						 "000100010101100111001100",
						 "000100010101100011100110",
						 "000100010110011001100000",
						 "000100010110010101111010",
						 "000100010110010010010100",
						 "000100010110001110101110",
						 "000100010110001011001000",
						 "000100010110000111100010",
						 "000100010110000011111100",
						 "000100010110000000010110",
						 "000100010101111100110000",
						 "000100010101111001001010",
						 "000100010101110101100100",
						 "000100010101110001111110",
						 "000100010101101110011000",
						 "000100010101101010110010",
						 "000100010101100111001100",
						 "000100010101100011100110",
						 "000100010110011001101111",
						 "000100010110010110001000",
						 "000100010110010010100001",
						 "000100010110001110111010",
						 "000100010110001011010011",
						 "000100010110000111101100",
						 "000100010110000100000101",
						 "000100010110000000011110",
						 "000100010101111100110111",
						 "000100010101111001010000",
						 "000100010101110101101001",
						 "000100010101110010000010",
						 "000100010101101110011011",
						 "000100010101101010110100",
						 "000100010101100111001101",
						 "000100010101100011100110",
						 "000100010011110110110001",
						 "000100010011110011001010",
						 "000100010011101111100011",
						 "000100010011101011111100",
						 "000100010011101000010101",
						 "000100010011100100101110",
						 "000100010011100001000111",
						 "000100010011011101100000",
						 "000100010011011001111001",
						 "000100010011010110010010",
						 "000100010011010010101011",
						 "000100010011001111000100",
						 "000100010011001011011101",
						 "000100010011000111110110",
						 "000100010011000100001111",
						 "000100010011000000101000",
						 "000100010011110110110001",
						 "000100010011110011001010",
						 "000100010011101111100011",
						 "000100010011101011111100",
						 "000100010011101000010101",
						 "000100010011100100101110",
						 "000100010011100001000111",
						 "000100010011011101100000",
						 "000100010011011001111001",
						 "000100010011010110010010",
						 "000100010011010010101011",
						 "000100010011001111000100",
						 "000100010011001011011101",
						 "000100010011000111110110",
						 "000100010011000100001111",
						 "000100010011000000101000",
						 "000100010011110110110001",
						 "000100010011110011001010",
						 "000100010011101111100011",
						 "000100010011101011111100",
						 "000100010011101000010101",
						 "000100010011100100101110",
						 "000100010011100001000111",
						 "000100010011011101100000",
						 "000100010011011001111001",
						 "000100010011010110010010",
						 "000100010011010010101011",
						 "000100010011001111000100",
						 "000100010011001011011101",
						 "000100010011000111110110",
						 "000100010011000100001111",
						 "000100010011000000101000",
						 "000100010001010011110011",
						 "000100010001010000001100",
						 "000100010001001100100101",
						 "000100010001001000111110",
						 "000100010001000101010111",
						 "000100010001000001110000",
						 "000100010000111110001001",
						 "000100010000111010100010",
						 "000100010000110110111011",
						 "000100010000110011010100",
						 "000100010000101111101101",
						 "000100010000101100000110",
						 "000100010000101000011111",
						 "000100010000100100111000",
						 "000100010000100001010001",
						 "000100010000011101101010",
						 "000100010001010011110011",
						 "000100010001010000001100",
						 "000100010001001100100101",
						 "000100010001001000111110",
						 "000100010001000101010111",
						 "000100010001000001110000",
						 "000100010000111110001001",
						 "000100010000111010100010",
						 "000100010000110110111011",
						 "000100010000110011010100",
						 "000100010000101111101101",
						 "000100010000101100000110",
						 "000100010000101000011111",
						 "000100010000100100111000",
						 "000100010000100001010001",
						 "000100010000011101101010",
						 "000100010001010100000010",
						 "000100010001010000011010",
						 "000100010001001100110010",
						 "000100010001001001001010",
						 "000100010001000101100010",
						 "000100010001000001111010",
						 "000100010000111110010010",
						 "000100010000111010101010",
						 "000100010000110111000010",
						 "000100010000110011011010",
						 "000100010000101111110010",
						 "000100010000101100001010",
						 "000100010000101000100010",
						 "000100010000100100111010",
						 "000100010000100001010010",
						 "000100010000011101101010",
						 "000100001110110001000100",
						 "000100001110101101011100",
						 "000100001110101001110100",
						 "000100001110100110001100",
						 "000100001110100010100100",
						 "000100001110011110111100",
						 "000100001110011011010100",
						 "000100001110010111101100",
						 "000100001110010100000100",
						 "000100001110010000011100",
						 "000100001110001100110100",
						 "000100001110001001001100",
						 "000100001110000101100100",
						 "000100001110000001111100",
						 "000100001101111110010100",
						 "000100001101111010101100",
						 "000100001110110001000100",
						 "000100001110101101011100",
						 "000100001110101001110100",
						 "000100001110100110001100",
						 "000100001110100010100100",
						 "000100001110011110111100",
						 "000100001110011011010100",
						 "000100001110010111101100",
						 "000100001110010100000100",
						 "000100001110010000011100",
						 "000100001110001100110100",
						 "000100001110001001001100",
						 "000100001110000101100100",
						 "000100001110000001111100",
						 "000100001101111110010100",
						 "000100001101111010101100",
						 "000100001100001110000110",
						 "000100001100001010011110",
						 "000100001100000110110110",
						 "000100001100000011001110",
						 "000100001011111111100110",
						 "000100001011111011111110",
						 "000100001011111000010110",
						 "000100001011110100101110",
						 "000100001011110001000110",
						 "000100001011101101011110",
						 "000100001011101001110110",
						 "000100001011100110001110",
						 "000100001011100010100110",
						 "000100001011011110111110",
						 "000100001011011011010110",
						 "000100001011010111101110",
						 "000100001100001110000110",
						 "000100001100001010011110",
						 "000100001100000110110110",
						 "000100001100000011001110",
						 "000100001011111111100110",
						 "000100001011111011111110",
						 "000100001011111000010110",
						 "000100001011110100101110",
						 "000100001011110001000110",
						 "000100001011101101011110",
						 "000100001011101001110110",
						 "000100001011100110001110",
						 "000100001011100010100110",
						 "000100001011011110111110",
						 "000100001011011011010110",
						 "000100001011010111101110",
						 "000100001100001110000110",
						 "000100001100001010011110",
						 "000100001100000110110110",
						 "000100001100000011001110",
						 "000100001011111111100110",
						 "000100001011111011111110",
						 "000100001011111000010110",
						 "000100001011110100101110",
						 "000100001011110001000110",
						 "000100001011101101011110",
						 "000100001011101001110110",
						 "000100001011100110001110",
						 "000100001011100010100110",
						 "000100001011011110111110",
						 "000100001011011011010110",
						 "000100001011010111101110",
						 "000100001001101011010111",
						 "000100001001100111101110",
						 "000100001001100100000101",
						 "000100001001100000011100",
						 "000100001001011100110011",
						 "000100001001011001001010",
						 "000100001001010101100001",
						 "000100001001010001111000",
						 "000100001001001110001111",
						 "000100001001001010100110",
						 "000100001001000110111101",
						 "000100001001000011010100",
						 "000100001000111111101011",
						 "000100001000111100000010",
						 "000100001000111000011001",
						 "000100001000110100110000",
						 "000100001001101011010111",
						 "000100001001100111101110",
						 "000100001001100100000101",
						 "000100001001100000011100",
						 "000100001001011100110011",
						 "000100001001011001001010",
						 "000100001001010101100001",
						 "000100001001010001111000",
						 "000100001001001110001111",
						 "000100001001001010100110",
						 "000100001001000110111101",
						 "000100001001000011010100",
						 "000100001000111111101011",
						 "000100001000111100000010",
						 "000100001000111000011001",
						 "000100001000110100110000",
						 "000100001001101011010111",
						 "000100001001100111101110",
						 "000100001001100100000101",
						 "000100001001100000011100",
						 "000100001001011100110011",
						 "000100001001011001001010",
						 "000100001001010101100001",
						 "000100001001010001111000",
						 "000100001001001110001111",
						 "000100001001001010100110",
						 "000100001001000110111101",
						 "000100001001000011010100",
						 "000100001000111111101011",
						 "000100001000111100000010",
						 "000100001000111000011001",
						 "000100001000110100110000",
						 "000100000111001000011001",
						 "000100000111000100110000",
						 "000100000111000001000111",
						 "000100000110111101011110",
						 "000100000110111001110101",
						 "000100000110110110001100",
						 "000100000110110010100011",
						 "000100000110101110111010",
						 "000100000110101011010001",
						 "000100000110100111101000",
						 "000100000110100011111111",
						 "000100000110100000010110",
						 "000100000110011100101101",
						 "000100000110011001000100",
						 "000100000110010101011011",
						 "000100000110010001110010",
						 "000100000111001000011001",
						 "000100000111000100110000",
						 "000100000111000001000111",
						 "000100000110111101011110",
						 "000100000110111001110101",
						 "000100000110110110001100",
						 "000100000110110010100011",
						 "000100000110101110111010",
						 "000100000110101011010001",
						 "000100000110100111101000",
						 "000100000110100011111111",
						 "000100000110100000010110",
						 "000100000110011100101101",
						 "000100000110011001000100",
						 "000100000110010101011011",
						 "000100000110010001110010",
						 "000100000111001000011001",
						 "000100000111000100110000",
						 "000100000111000001000111",
						 "000100000110111101011110",
						 "000100000110111001110101",
						 "000100000110110110001100",
						 "000100000110110010100011",
						 "000100000110101110111010",
						 "000100000110101011010001",
						 "000100000110100111101000",
						 "000100000110100011111111",
						 "000100000110100000010110",
						 "000100000110011100101101",
						 "000100000110011001000100",
						 "000100000110010101011011",
						 "000100000110010001110010",
						 "000100000100100101101010",
						 "000100000100100010000000",
						 "000100000100011110010110",
						 "000100000100011010101100",
						 "000100000100010111000010",
						 "000100000100010011011000",
						 "000100000100001111101110",
						 "000100000100001100000100",
						 "000100000100001000011010",
						 "000100000100000100110000",
						 "000100000100000001000110",
						 "000100000011111101011100",
						 "000100000011111001110010",
						 "000100000011110110001000",
						 "000100000011110010011110",
						 "000100000011101110110100",
						 "000100000100100101101010",
						 "000100000100100010000000",
						 "000100000100011110010110",
						 "000100000100011010101100",
						 "000100000100010111000010",
						 "000100000100010011011000",
						 "000100000100001111101110",
						 "000100000100001100000100",
						 "000100000100001000011010",
						 "000100000100000100110000",
						 "000100000100000001000110",
						 "000100000011111101011100",
						 "000100000011111001110010",
						 "000100000011110110001000",
						 "000100000011110010011110",
						 "000100000011101110110100",
						 "000100000100100101101010",
						 "000100000100100010000000",
						 "000100000100011110010110",
						 "000100000100011010101100",
						 "000100000100010111000010",
						 "000100000100010011011000",
						 "000100000100001111101110",
						 "000100000100001100000100",
						 "000100000100001000011010",
						 "000100000100000100110000",
						 "000100000100000001000110",
						 "000100000011111101011100",
						 "000100000011111001110010",
						 "000100000011110110001000",
						 "000100000011110010011110",
						 "000100000011101110110100",
						 "000100000010000010101100",
						 "000100000001111111000010",
						 "000100000001111011011000",
						 "000100000001110111101110",
						 "000100000001110100000100",
						 "000100000001110000011010",
						 "000100000001101100110000",
						 "000100000001101001000110",
						 "000100000001100101011100",
						 "000100000001100001110010",
						 "000100000001011110001000",
						 "000100000001011010011110",
						 "000100000001010110110100",
						 "000100000001010011001010",
						 "000100000001001111100000",
						 "000100000001001011110110",
						 "000100000010000010101100",
						 "000100000001111111000010",
						 "000100000001111011011000",
						 "000100000001110111101110",
						 "000100000001110100000100",
						 "000100000001110000011010",
						 "000100000001101100110000",
						 "000100000001101001000110",
						 "000100000001100101011100",
						 "000100000001100001110010",
						 "000100000001011110001000",
						 "000100000001011010011110",
						 "000100000001010110110100",
						 "000100000001010011001010",
						 "000100000001001111100000",
						 "000100000001001011110110",
						 "000011111111011111101110",
						 "000011111111011100000100",
						 "000011111111011000011010",
						 "000011111111010100110000",
						 "000011111111010001000110",
						 "000011111111001101011100",
						 "000011111111001001110010",
						 "000011111111000110001000",
						 "000011111111000010011110",
						 "000011111110111110110100",
						 "000011111110111011001010",
						 "000011111110110111100000",
						 "000011111110110011110110",
						 "000011111110110000001100",
						 "000011111110101100100010",
						 "000011111110101000111000",
						 "000011111111011111101110",
						 "000011111111011100000100",
						 "000011111111011000011010",
						 "000011111111010100110000",
						 "000011111111010001000110",
						 "000011111111001101011100",
						 "000011111111001001110010",
						 "000011111111000110001000",
						 "000011111111000010011110",
						 "000011111110111110110100",
						 "000011111110111011001010",
						 "000011111110110111100000",
						 "000011111110110011110110",
						 "000011111110110000001100",
						 "000011111110101100100010",
						 "000011111110101000111000",
						 "000011111111011111111101",
						 "000011111111011100010010",
						 "000011111111011000100111",
						 "000011111111010100111100",
						 "000011111111010001010001",
						 "000011111111001101100110",
						 "000011111111001001111011",
						 "000011111111000110010000",
						 "000011111111000010100101",
						 "000011111110111110111010",
						 "000011111110111011001111",
						 "000011111110110111100100",
						 "000011111110110011111001",
						 "000011111110110000001110",
						 "000011111110101100100011",
						 "000011111110101000111000",
						 "000011111100111100111111",
						 "000011111100111001010100",
						 "000011111100110101101001",
						 "000011111100110001111110",
						 "000011111100101110010011",
						 "000011111100101010101000",
						 "000011111100100110111101",
						 "000011111100100011010010",
						 "000011111100011111100111",
						 "000011111100011011111100",
						 "000011111100011000010001",
						 "000011111100010100100110",
						 "000011111100010000111011",
						 "000011111100001101010000",
						 "000011111100001001100101",
						 "000011111100000101111010",
						 "000011111100111100111111",
						 "000011111100111001010100",
						 "000011111100110101101001",
						 "000011111100110001111110",
						 "000011111100101110010011",
						 "000011111100101010101000",
						 "000011111100100110111101",
						 "000011111100100011010010",
						 "000011111100011111100111",
						 "000011111100011011111100",
						 "000011111100011000010001",
						 "000011111100010100100110",
						 "000011111100010000111011",
						 "000011111100001101010000",
						 "000011111100001001100101",
						 "000011111100000101111010",
						 "000011111100111100111111",
						 "000011111100111001010100",
						 "000011111100110101101001",
						 "000011111100110001111110",
						 "000011111100101110010011",
						 "000011111100101010101000",
						 "000011111100100110111101",
						 "000011111100100011010010",
						 "000011111100011111100111",
						 "000011111100011011111100",
						 "000011111100011000010001",
						 "000011111100010100100110",
						 "000011111100010000111011",
						 "000011111100001101010000",
						 "000011111100001001100101",
						 "000011111100000101111010",
						 "000011111010011010000001",
						 "000011111010010110010110",
						 "000011111010010010101011",
						 "000011111010001111000000",
						 "000011111010001011010101",
						 "000011111010000111101010",
						 "000011111010000011111111",
						 "000011111010000000010100",
						 "000011111001111100101001",
						 "000011111001111000111110",
						 "000011111001110101010011",
						 "000011111001110001101000",
						 "000011111001101101111101",
						 "000011111001101010010010",
						 "000011111001100110100111",
						 "000011111001100010111100",
						 "000011111010011010000001",
						 "000011111010010110010110",
						 "000011111010010010101011",
						 "000011111010001111000000",
						 "000011111010001011010101",
						 "000011111010000111101010",
						 "000011111010000011111111",
						 "000011111010000000010100",
						 "000011111001111100101001",
						 "000011111001111000111110",
						 "000011111001110101010011",
						 "000011111001110001101000",
						 "000011111001101101111101",
						 "000011111001101010010010",
						 "000011111001100110100111",
						 "000011111001100010111100",
						 "000011111010011010010000",
						 "000011111010010110100100",
						 "000011111010010010111000",
						 "000011111010001111001100",
						 "000011111010001011100000",
						 "000011111010000111110100",
						 "000011111010000100001000",
						 "000011111010000000011100",
						 "000011111001111100110000",
						 "000011111001111001000100",
						 "000011111001110101011000",
						 "000011111001110001101100",
						 "000011111001101110000000",
						 "000011111001101010010100",
						 "000011111001100110101000",
						 "000011111001100010111100",
						 "000011110111110111010010",
						 "000011110111110011100110",
						 "000011110111101111111010",
						 "000011110111101100001110",
						 "000011110111101000100010",
						 "000011110111100100110110",
						 "000011110111100001001010",
						 "000011110111011101011110",
						 "000011110111011001110010",
						 "000011110111010110000110",
						 "000011110111010010011010",
						 "000011110111001110101110",
						 "000011110111001011000010",
						 "000011110111000111010110",
						 "000011110111000011101010",
						 "000011110110111111111110",
						 "000011110111110111010010",
						 "000011110111110011100110",
						 "000011110111101111111010",
						 "000011110111101100001110",
						 "000011110111101000100010",
						 "000011110111100100110110",
						 "000011110111100001001010",
						 "000011110111011101011110",
						 "000011110111011001110010",
						 "000011110111010110000110",
						 "000011110111010010011010",
						 "000011110111001110101110",
						 "000011110111001011000010",
						 "000011110111000111010110",
						 "000011110111000011101010",
						 "000011110110111111111110",
						 "000011110111110111010010",
						 "000011110111110011100110",
						 "000011110111101111111010",
						 "000011110111101100001110",
						 "000011110111101000100010",
						 "000011110111100100110110",
						 "000011110111100001001010",
						 "000011110111011101011110",
						 "000011110111011001110010",
						 "000011110111010110000110",
						 "000011110111010010011010",
						 "000011110111001110101110",
						 "000011110111001011000010",
						 "000011110111000111010110",
						 "000011110111000011101010",
						 "000011110110111111111110",
						 "000011110101010100010100",
						 "000011110101010000101000",
						 "000011110101001100111100",
						 "000011110101001001010000",
						 "000011110101000101100100",
						 "000011110101000001111000",
						 "000011110100111110001100",
						 "000011110100111010100000",
						 "000011110100110110110100",
						 "000011110100110011001000",
						 "000011110100101111011100",
						 "000011110100101011110000",
						 "000011110100101000000100",
						 "000011110100100100011000",
						 "000011110100100000101100",
						 "000011110100011101000000",
						 "000011110101010100010100",
						 "000011110101010000101000",
						 "000011110101001100111100",
						 "000011110101001001010000",
						 "000011110101000101100100",
						 "000011110101000001111000",
						 "000011110100111110001100",
						 "000011110100111010100000",
						 "000011110100110110110100",
						 "000011110100110011001000",
						 "000011110100101111011100",
						 "000011110100101011110000",
						 "000011110100101000000100",
						 "000011110100100100011000",
						 "000011110100100000101100",
						 "000011110100011101000000",
						 "000011110010110001010110",
						 "000011110010101101101010",
						 "000011110010101001111110",
						 "000011110010100110010010",
						 "000011110010100010100110",
						 "000011110010011110111010",
						 "000011110010011011001110",
						 "000011110010010111100010",
						 "000011110010010011110110",
						 "000011110010010000001010",
						 "000011110010001100011110",
						 "000011110010001000110010",
						 "000011110010000101000110",
						 "000011110010000001011010",
						 "000011110001111101101110",
						 "000011110001111010000010",
						 "000011110010110001100101",
						 "000011110010101101111000",
						 "000011110010101010001011",
						 "000011110010100110011110",
						 "000011110010100010110001",
						 "000011110010011111000100",
						 "000011110010011011010111",
						 "000011110010010111101010",
						 "000011110010010011111101",
						 "000011110010010000010000",
						 "000011110010001100100011",
						 "000011110010001000110110",
						 "000011110010000101001001",
						 "000011110010000001011100",
						 "000011110001111101101111",
						 "000011110001111010000010",
						 "000011110010110001100101",
						 "000011110010101101111000",
						 "000011110010101010001011",
						 "000011110010100110011110",
						 "000011110010100010110001",
						 "000011110010011111000100",
						 "000011110010011011010111",
						 "000011110010010111101010",
						 "000011110010010011111101",
						 "000011110010010000010000",
						 "000011110010001100100011",
						 "000011110010001000110110",
						 "000011110010000101001001",
						 "000011110010000001011100",
						 "000011110001111101101111",
						 "000011110001111010000010",
						 "000011110000001110100111",
						 "000011110000001010111010",
						 "000011110000000111001101",
						 "000011110000000011100000",
						 "000011101111111111110011",
						 "000011101111111100000110",
						 "000011101111111000011001",
						 "000011101111110100101100",
						 "000011101111110000111111",
						 "000011101111101101010010",
						 "000011101111101001100101",
						 "000011101111100101111000",
						 "000011101111100010001011",
						 "000011101111011110011110",
						 "000011101111011010110001",
						 "000011101111010111000100",
						 "000011110000001110100111",
						 "000011110000001010111010",
						 "000011110000000111001101",
						 "000011110000000011100000",
						 "000011101111111111110011",
						 "000011101111111100000110",
						 "000011101111111000011001",
						 "000011101111110100101100",
						 "000011101111110000111111",
						 "000011101111101101010010",
						 "000011101111101001100101",
						 "000011101111100101111000",
						 "000011101111100010001011",
						 "000011101111011110011110",
						 "000011101111011010110001",
						 "000011101111010111000100",
						 "000011110000001110100111",
						 "000011110000001010111010",
						 "000011110000000111001101",
						 "000011110000000011100000",
						 "000011101111111111110011",
						 "000011101111111100000110",
						 "000011101111111000011001",
						 "000011101111110100101100",
						 "000011101111110000111111",
						 "000011101111101101010010",
						 "000011101111101001100101",
						 "000011101111100101111000",
						 "000011101111100010001011",
						 "000011101111011110011110",
						 "000011101111011010110001",
						 "000011101111010111000100",
						 "000011101101101011101001",
						 "000011101101100111111100",
						 "000011101101100100001111",
						 "000011101101100000100010",
						 "000011101101011100110101",
						 "000011101101011001001000",
						 "000011101101010101011011",
						 "000011101101010001101110",
						 "000011101101001110000001",
						 "000011101101001010010100",
						 "000011101101000110100111",
						 "000011101101000010111010",
						 "000011101100111111001101",
						 "000011101100111011100000",
						 "000011101100110111110011",
						 "000011101100110100000110",
						 "000011101101101011101001",
						 "000011101101100111111100",
						 "000011101101100100001111",
						 "000011101101100000100010",
						 "000011101101011100110101",
						 "000011101101011001001000",
						 "000011101101010101011011",
						 "000011101101010001101110",
						 "000011101101001110000001",
						 "000011101101001010010100",
						 "000011101101000110100111",
						 "000011101101000010111010",
						 "000011101100111111001101",
						 "000011101100111011100000",
						 "000011101100110111110011",
						 "000011101100110100000110",
						 "000011101101101011111000",
						 "000011101101101000001010",
						 "000011101101100100011100",
						 "000011101101100000101110",
						 "000011101101011101000000",
						 "000011101101011001010010",
						 "000011101101010101100100",
						 "000011101101010001110110",
						 "000011101101001110001000",
						 "000011101101001010011010",
						 "000011101101000110101100",
						 "000011101101000010111110",
						 "000011101100111111010000",
						 "000011101100111011100010",
						 "000011101100110111110100",
						 "000011101100110100000110",
						 "000011101011001000111010",
						 "000011101011000101001100",
						 "000011101011000001011110",
						 "000011101010111101110000",
						 "000011101010111010000010",
						 "000011101010110110010100",
						 "000011101010110010100110",
						 "000011101010101110111000",
						 "000011101010101011001010",
						 "000011101010100111011100",
						 "000011101010100011101110",
						 "000011101010100000000000",
						 "000011101010011100010010",
						 "000011101010011000100100",
						 "000011101010010100110110",
						 "000011101010010001001000",
						 "000011101011001000111010",
						 "000011101011000101001100",
						 "000011101011000001011110",
						 "000011101010111101110000",
						 "000011101010111010000010",
						 "000011101010110110010100",
						 "000011101010110010100110",
						 "000011101010101110111000",
						 "000011101010101011001010",
						 "000011101010100111011100",
						 "000011101010100011101110",
						 "000011101010100000000000",
						 "000011101010011100010010",
						 "000011101010011000100100",
						 "000011101010010100110110",
						 "000011101010010001001000",
						 "000011101000100101111100",
						 "000011101000100010001110",
						 "000011101000011110100000",
						 "000011101000011010110010",
						 "000011101000010111000100",
						 "000011101000010011010110",
						 "000011101000001111101000",
						 "000011101000001011111010",
						 "000011101000001000001100",
						 "000011101000000100011110",
						 "000011101000000000110000",
						 "000011100111111101000010",
						 "000011100111111001010100",
						 "000011100111110101100110",
						 "000011100111110001111000",
						 "000011100111101110001010",
						 "000011101000100101111100",
						 "000011101000100010001110",
						 "000011101000011110100000",
						 "000011101000011010110010",
						 "000011101000010111000100",
						 "000011101000010011010110",
						 "000011101000001111101000",
						 "000011101000001011111010",
						 "000011101000001000001100",
						 "000011101000000100011110",
						 "000011101000000000110000",
						 "000011100111111101000010",
						 "000011100111111001010100",
						 "000011100111110101100110",
						 "000011100111110001111000",
						 "000011100111101110001010",
						 "000011101000100101111100",
						 "000011101000100010001110",
						 "000011101000011110100000",
						 "000011101000011010110010",
						 "000011101000010111000100",
						 "000011101000010011010110",
						 "000011101000001111101000",
						 "000011101000001011111010",
						 "000011101000001000001100",
						 "000011101000000100011110",
						 "000011101000000000110000",
						 "000011100111111101000010",
						 "000011100111111001010100",
						 "000011100111110101100110",
						 "000011100111110001111000",
						 "000011100111101110001010",
						 "000011100110000010111110",
						 "000011100101111111010000",
						 "000011100101111011100010",
						 "000011100101110111110100",
						 "000011100101110100000110",
						 "000011100101110000011000",
						 "000011100101101100101010",
						 "000011100101101000111100",
						 "000011100101100101001110",
						 "000011100101100001100000",
						 "000011100101011101110010",
						 "000011100101011010000100",
						 "000011100101010110010110",
						 "000011100101010010101000",
						 "000011100101001110111010",
						 "000011100101001011001100",
						 "000011100110000011001101",
						 "000011100101111111011110",
						 "000011100101111011101111",
						 "000011100101111000000000",
						 "000011100101110100010001",
						 "000011100101110000100010",
						 "000011100101101100110011",
						 "000011100101101001000100",
						 "000011100101100101010101",
						 "000011100101100001100110",
						 "000011100101011101110111",
						 "000011100101011010001000",
						 "000011100101010110011001",
						 "000011100101010010101010",
						 "000011100101001110111011",
						 "000011100101001011001100",
						 "000011100110000011001101",
						 "000011100101111111011110",
						 "000011100101111011101111",
						 "000011100101111000000000",
						 "000011100101110100010001",
						 "000011100101110000100010",
						 "000011100101101100110011",
						 "000011100101101001000100",
						 "000011100101100101010101",
						 "000011100101100001100110",
						 "000011100101011101110111",
						 "000011100101011010001000",
						 "000011100101010110011001",
						 "000011100101010010101010",
						 "000011100101001110111011",
						 "000011100101001011001100",
						 "000011100011100000001111",
						 "000011100011011100100000",
						 "000011100011011000110001",
						 "000011100011010101000010",
						 "000011100011010001010011",
						 "000011100011001101100100",
						 "000011100011001001110101",
						 "000011100011000110000110",
						 "000011100011000010010111",
						 "000011100010111110101000",
						 "000011100010111010111001",
						 "000011100010110111001010",
						 "000011100010110011011011",
						 "000011100010101111101100",
						 "000011100010101011111101",
						 "000011100010101000001110",
						 "000011100011100000001111",
						 "000011100011011100100000",
						 "000011100011011000110001",
						 "000011100011010101000010",
						 "000011100011010001010011",
						 "000011100011001101100100",
						 "000011100011001001110101",
						 "000011100011000110000110",
						 "000011100011000010010111",
						 "000011100010111110101000",
						 "000011100010111010111001",
						 "000011100010110111001010",
						 "000011100010110011011011",
						 "000011100010101111101100",
						 "000011100010101011111101",
						 "000011100010101000001110",
						 "000011100000111101010001",
						 "000011100000111001100010",
						 "000011100000110101110011",
						 "000011100000110010000100",
						 "000011100000101110010101",
						 "000011100000101010100110",
						 "000011100000100110110111",
						 "000011100000100011001000",
						 "000011100000011111011001",
						 "000011100000011011101010",
						 "000011100000010111111011",
						 "000011100000010100001100",
						 "000011100000010000011101",
						 "000011100000001100101110",
						 "000011100000001000111111",
						 "000011100000000101010000",
						 "000011100000111101010001",
						 "000011100000111001100010",
						 "000011100000110101110011",
						 "000011100000110010000100",
						 "000011100000101110010101",
						 "000011100000101010100110",
						 "000011100000100110110111",
						 "000011100000100011001000",
						 "000011100000011111011001",
						 "000011100000011011101010",
						 "000011100000010111111011",
						 "000011100000010100001100",
						 "000011100000010000011101",
						 "000011100000001100101110",
						 "000011100000001000111111",
						 "000011100000000101010000",
						 "000011100000111101010001",
						 "000011100000111001100010",
						 "000011100000110101110011",
						 "000011100000110010000100",
						 "000011100000101110010101",
						 "000011100000101010100110",
						 "000011100000100110110111",
						 "000011100000100011001000",
						 "000011100000011111011001",
						 "000011100000011011101010",
						 "000011100000010111111011",
						 "000011100000010100001100",
						 "000011100000010000011101",
						 "000011100000001100101110",
						 "000011100000001000111111",
						 "000011100000000101010000",
						 "000011011110011010010011",
						 "000011011110010110100100",
						 "000011011110010010110101",
						 "000011011110001111000110",
						 "000011011110001011010111",
						 "000011011110000111101000",
						 "000011011110000011111001",
						 "000011011110000000001010",
						 "000011011101111100011011",
						 "000011011101111000101100",
						 "000011011101110100111101",
						 "000011011101110001001110",
						 "000011011101101101011111",
						 "000011011101101001110000",
						 "000011011101100110000001",
						 "000011011101100010010010",
						 "000011011110011010100010",
						 "000011011110010110110010",
						 "000011011110010011000010",
						 "000011011110001111010010",
						 "000011011110001011100010",
						 "000011011110000111110010",
						 "000011011110000100000010",
						 "000011011110000000010010",
						 "000011011101111100100010",
						 "000011011101111000110010",
						 "000011011101110101000010",
						 "000011011101110001010010",
						 "000011011101101101100010",
						 "000011011101101001110010",
						 "000011011101100110000010",
						 "000011011101100010010010",
						 "000011011110011010100010",
						 "000011011110010110110010",
						 "000011011110010011000010",
						 "000011011110001111010010",
						 "000011011110001011100010",
						 "000011011110000111110010",
						 "000011011110000100000010",
						 "000011011110000000010010",
						 "000011011101111100100010",
						 "000011011101111000110010",
						 "000011011101110101000010",
						 "000011011101110001010010",
						 "000011011101101101100010",
						 "000011011101101001110010",
						 "000011011101100110000010",
						 "000011011101100010010010",
						 "000011011011110111100100",
						 "000011011011110011110100",
						 "000011011011110000000100",
						 "000011011011101100010100",
						 "000011011011101000100100",
						 "000011011011100100110100",
						 "000011011011100001000100",
						 "000011011011011101010100",
						 "000011011011011001100100",
						 "000011011011010101110100",
						 "000011011011010010000100",
						 "000011011011001110010100",
						 "000011011011001010100100",
						 "000011011011000110110100",
						 "000011011011000011000100",
						 "000011011010111111010100",
						 "000011011011110111100100",
						 "000011011011110011110100",
						 "000011011011110000000100",
						 "000011011011101100010100",
						 "000011011011101000100100",
						 "000011011011100100110100",
						 "000011011011100001000100",
						 "000011011011011101010100",
						 "000011011011011001100100",
						 "000011011011010101110100",
						 "000011011011010010000100",
						 "000011011011001110010100",
						 "000011011011001010100100",
						 "000011011011000110110100",
						 "000011011011000011000100",
						 "000011011010111111010100",
						 "000011011011110111100100",
						 "000011011011110011110100",
						 "000011011011110000000100",
						 "000011011011101100010100",
						 "000011011011101000100100",
						 "000011011011100100110100",
						 "000011011011100001000100",
						 "000011011011011101010100",
						 "000011011011011001100100",
						 "000011011011010101110100",
						 "000011011011010010000100",
						 "000011011011001110010100",
						 "000011011011001010100100",
						 "000011011011000110110100",
						 "000011011011000011000100",
						 "000011011010111111010100",
						 "000011011001010100100110",
						 "000011011001010000110110",
						 "000011011001001101000110",
						 "000011011001001001010110",
						 "000011011001000101100110",
						 "000011011001000001110110",
						 "000011011000111110000110",
						 "000011011000111010010110",
						 "000011011000110110100110",
						 "000011011000110010110110",
						 "000011011000101111000110",
						 "000011011000101011010110",
						 "000011011000100111100110",
						 "000011011000100011110110",
						 "000011011000100000000110",
						 "000011011000011100010110",
						 "000011011001010100100110",
						 "000011011001010000110110",
						 "000011011001001101000110",
						 "000011011001001001010110",
						 "000011011001000101100110",
						 "000011011001000001110110",
						 "000011011000111110000110",
						 "000011011000111010010110",
						 "000011011000110110100110",
						 "000011011000110010110110",
						 "000011011000101111000110",
						 "000011011000101011010110",
						 "000011011000100111100110",
						 "000011011000100011110110",
						 "000011011000100000000110",
						 "000011011000011100010110",
						 "000011010110110001110111",
						 "000011010110101110000110",
						 "000011010110101010010101",
						 "000011010110100110100100",
						 "000011010110100010110011",
						 "000011010110011111000010",
						 "000011010110011011010001",
						 "000011010110010111100000",
						 "000011010110010011101111",
						 "000011010110001111111110",
						 "000011010110001100001101",
						 "000011010110001000011100",
						 "000011010110000100101011",
						 "000011010110000000111010",
						 "000011010101111101001001",
						 "000011010101111001011000",
						 "000011010110110001110111",
						 "000011010110101110000110",
						 "000011010110101010010101",
						 "000011010110100110100100",
						 "000011010110100010110011",
						 "000011010110011111000010",
						 "000011010110011011010001",
						 "000011010110010111100000",
						 "000011010110010011101111",
						 "000011010110001111111110",
						 "000011010110001100001101",
						 "000011010110001000011100",
						 "000011010110000100101011",
						 "000011010110000000111010",
						 "000011010101111101001001",
						 "000011010101111001011000",
						 "000011010110110001110111",
						 "000011010110101110000110",
						 "000011010110101010010101",
						 "000011010110100110100100",
						 "000011010110100010110011",
						 "000011010110011111000010",
						 "000011010110011011010001",
						 "000011010110010111100000",
						 "000011010110010011101111",
						 "000011010110001111111110",
						 "000011010110001100001101",
						 "000011010110001000011100",
						 "000011010110000100101011",
						 "000011010110000000111010",
						 "000011010101111101001001",
						 "000011010101111001011000",
						 "000011010100001110111001",
						 "000011010100001011001000",
						 "000011010100000111010111",
						 "000011010100000011100110",
						 "000011010011111111110101",
						 "000011010011111100000100",
						 "000011010011111000010011",
						 "000011010011110100100010",
						 "000011010011110000110001",
						 "000011010011101101000000",
						 "000011010011101001001111",
						 "000011010011100101011110",
						 "000011010011100001101101",
						 "000011010011011101111100",
						 "000011010011011010001011",
						 "000011010011010110011010",
						 "000011010100001110111001",
						 "000011010100001011001000",
						 "000011010100000111010111",
						 "000011010100000011100110",
						 "000011010011111111110101",
						 "000011010011111100000100",
						 "000011010011111000010011",
						 "000011010011110100100010",
						 "000011010011110000110001",
						 "000011010011101101000000",
						 "000011010011101001001111",
						 "000011010011100101011110",
						 "000011010011100001101101",
						 "000011010011011101111100",
						 "000011010011011010001011",
						 "000011010011010110011010",
						 "000011010100001110111001",
						 "000011010100001011001000",
						 "000011010100000111010111",
						 "000011010100000011100110",
						 "000011010011111111110101",
						 "000011010011111100000100",
						 "000011010011111000010011",
						 "000011010011110100100010",
						 "000011010011110000110001",
						 "000011010011101101000000",
						 "000011010011101001001111",
						 "000011010011100101011110",
						 "000011010011100001101101",
						 "000011010011011101111100",
						 "000011010011011010001011",
						 "000011010011010110011010",
						 "000011010001101011111011",
						 "000011010001101000001010",
						 "000011010001100100011001",
						 "000011010001100000101000",
						 "000011010001011100110111",
						 "000011010001011001000110",
						 "000011010001010101010101",
						 "000011010001010001100100",
						 "000011010001001101110011",
						 "000011010001001010000010",
						 "000011010001000110010001",
						 "000011010001000010100000",
						 "000011010000111110101111",
						 "000011010000111010111110",
						 "000011010000110111001101",
						 "000011010000110011011100",
						 "000011010001101011111011",
						 "000011010001101000001010",
						 "000011010001100100011001",
						 "000011010001100000101000",
						 "000011010001011100110111",
						 "000011010001011001000110",
						 "000011010001010101010101",
						 "000011010001010001100100",
						 "000011010001001101110011",
						 "000011010001001010000010",
						 "000011010001000110010001",
						 "000011010001000010100000",
						 "000011010000111110101111",
						 "000011010000111010111110",
						 "000011010000110111001101",
						 "000011010000110011011100",
						 "000011001111001001001100",
						 "000011001111000101011010",
						 "000011001111000001101000",
						 "000011001110111101110110",
						 "000011001110111010000100",
						 "000011001110110110010010",
						 "000011001110110010100000",
						 "000011001110101110101110",
						 "000011001110101010111100",
						 "000011001110100111001010",
						 "000011001110100011011000",
						 "000011001110011111100110",
						 "000011001110011011110100",
						 "000011001110011000000010",
						 "000011001110010100010000",
						 "000011001110010000011110",
						 "000011001111001001001100",
						 "000011001111000101011010",
						 "000011001111000001101000",
						 "000011001110111101110110",
						 "000011001110111010000100",
						 "000011001110110110010010",
						 "000011001110110010100000",
						 "000011001110101110101110",
						 "000011001110101010111100",
						 "000011001110100111001010",
						 "000011001110100011011000",
						 "000011001110011111100110",
						 "000011001110011011110100",
						 "000011001110011000000010",
						 "000011001110010100010000",
						 "000011001110010000011110",
						 "000011001111001001001100",
						 "000011001111000101011010",
						 "000011001111000001101000",
						 "000011001110111101110110",
						 "000011001110111010000100",
						 "000011001110110110010010",
						 "000011001110110010100000",
						 "000011001110101110101110",
						 "000011001110101010111100",
						 "000011001110100111001010",
						 "000011001110100011011000",
						 "000011001110011111100110",
						 "000011001110011011110100",
						 "000011001110011000000010",
						 "000011001110010100010000",
						 "000011001110010000011110",
						 "000011001100100110001110",
						 "000011001100100010011100",
						 "000011001100011110101010",
						 "000011001100011010111000",
						 "000011001100010111000110",
						 "000011001100010011010100",
						 "000011001100001111100010",
						 "000011001100001011110000",
						 "000011001100000111111110",
						 "000011001100000100001100",
						 "000011001100000000011010",
						 "000011001011111100101000",
						 "000011001011111000110110",
						 "000011001011110101000100",
						 "000011001011110001010010",
						 "000011001011101101100000",
						 "000011001100100110001110",
						 "000011001100100010011100",
						 "000011001100011110101010",
						 "000011001100011010111000",
						 "000011001100010111000110",
						 "000011001100010011010100",
						 "000011001100001111100010",
						 "000011001100001011110000",
						 "000011001100000111111110",
						 "000011001100000100001100",
						 "000011001100000000011010",
						 "000011001011111100101000",
						 "000011001011111000110110",
						 "000011001011110101000100",
						 "000011001011110001010010",
						 "000011001011101101100000",
						 "000011001100100110001110",
						 "000011001100100010011100",
						 "000011001100011110101010",
						 "000011001100011010111000",
						 "000011001100010111000110",
						 "000011001100010011010100",
						 "000011001100001111100010",
						 "000011001100001011110000",
						 "000011001100000111111110",
						 "000011001100000100001100",
						 "000011001100000000011010",
						 "000011001011111100101000",
						 "000011001011111000110110",
						 "000011001011110101000100",
						 "000011001011110001010010",
						 "000011001011101101100000",
						 "000011001010000011010000",
						 "000011001001111111011110",
						 "000011001001111011101100",
						 "000011001001110111111010",
						 "000011001001110100001000",
						 "000011001001110000010110",
						 "000011001001101100100100",
						 "000011001001101000110010",
						 "000011001001100101000000",
						 "000011001001100001001110",
						 "000011001001011101011100",
						 "000011001001011001101010",
						 "000011001001010101111000",
						 "000011001001010010000110",
						 "000011001001001110010100",
						 "000011001001001010100010",
						 "000011001010000011010000",
						 "000011001001111111011110",
						 "000011001001111011101100",
						 "000011001001110111111010",
						 "000011001001110100001000",
						 "000011001001110000010110",
						 "000011001001101100100100",
						 "000011001001101000110010",
						 "000011001001100101000000",
						 "000011001001100001001110",
						 "000011001001011101011100",
						 "000011001001011001101010",
						 "000011001001010101111000",
						 "000011001001010010000110",
						 "000011001001001110010100",
						 "000011001001001010100010",
						 "000011001010000011011111",
						 "000011001001111111101100",
						 "000011001001111011111001",
						 "000011001001111000000110",
						 "000011001001110100010011",
						 "000011001001110000100000",
						 "000011001001101100101101",
						 "000011001001101000111010",
						 "000011001001100101000111",
						 "000011001001100001010100",
						 "000011001001011101100001",
						 "000011001001011001101110",
						 "000011001001010101111011",
						 "000011001001010010001000",
						 "000011001001001110010101",
						 "000011001001001010100010",
						 "000011000111100000100001",
						 "000011000111011100101110",
						 "000011000111011000111011",
						 "000011000111010101001000",
						 "000011000111010001010101",
						 "000011000111001101100010",
						 "000011000111001001101111",
						 "000011000111000101111100",
						 "000011000111000010001001",
						 "000011000110111110010110",
						 "000011000110111010100011",
						 "000011000110110110110000",
						 "000011000110110010111101",
						 "000011000110101111001010",
						 "000011000110101011010111",
						 "000011000110100111100100",
						 "000011000111100000100001",
						 "000011000111011100101110",
						 "000011000111011000111011",
						 "000011000111010101001000",
						 "000011000111010001010101",
						 "000011000111001101100010",
						 "000011000111001001101111",
						 "000011000111000101111100",
						 "000011000111000010001001",
						 "000011000110111110010110",
						 "000011000110111010100011",
						 "000011000110110110110000",
						 "000011000110110010111101",
						 "000011000110101111001010",
						 "000011000110101011010111",
						 "000011000110100111100100",
						 "000011000100111101100011",
						 "000011000100111001110000",
						 "000011000100110101111101",
						 "000011000100110010001010",
						 "000011000100101110010111",
						 "000011000100101010100100",
						 "000011000100100110110001",
						 "000011000100100010111110",
						 "000011000100011111001011",
						 "000011000100011011011000",
						 "000011000100010111100101",
						 "000011000100010011110010",
						 "000011000100001111111111",
						 "000011000100001100001100",
						 "000011000100001000011001",
						 "000011000100000100100110",
						 "000011000100111101100011",
						 "000011000100111001110000",
						 "000011000100110101111101",
						 "000011000100110010001010",
						 "000011000100101110010111",
						 "000011000100101010100100",
						 "000011000100100110110001",
						 "000011000100100010111110",
						 "000011000100011111001011",
						 "000011000100011011011000",
						 "000011000100010111100101",
						 "000011000100010011110010",
						 "000011000100001111111111",
						 "000011000100001100001100",
						 "000011000100001000011001",
						 "000011000100000100100110",
						 "000011000100111101100011",
						 "000011000100111001110000",
						 "000011000100110101111101",
						 "000011000100110010001010",
						 "000011000100101110010111",
						 "000011000100101010100100",
						 "000011000100100110110001",
						 "000011000100100010111110",
						 "000011000100011111001011",
						 "000011000100011011011000",
						 "000011000100010111100101",
						 "000011000100010011110010",
						 "000011000100001111111111",
						 "000011000100001100001100",
						 "000011000100001000011001",
						 "000011000100000100100110",
						 "000011000010011010100101",
						 "000011000010010110110010",
						 "000011000010010010111111",
						 "000011000010001111001100",
						 "000011000010001011011001",
						 "000011000010000111100110",
						 "000011000010000011110011",
						 "000011000010000000000000",
						 "000011000001111100001101",
						 "000011000001111000011010",
						 "000011000001110100100111",
						 "000011000001110000110100",
						 "000011000001101101000001",
						 "000011000001101001001110",
						 "000011000001100101011011",
						 "000011000001100001101000",
						 "000011000010011010100101",
						 "000011000010010110110010",
						 "000011000010010010111111",
						 "000011000010001111001100",
						 "000011000010001011011001",
						 "000011000010000111100110",
						 "000011000010000011110011",
						 "000011000010000000000000",
						 "000011000001111100001101",
						 "000011000001111000011010",
						 "000011000001110100100111",
						 "000011000001110000110100",
						 "000011000001101101000001",
						 "000011000001101001001110",
						 "000011000001100101011011",
						 "000011000001100001101000",
						 "000011000010011010110100",
						 "000011000010010111000000",
						 "000011000010010011001100",
						 "000011000010001111011000",
						 "000011000010001011100100",
						 "000011000010000111110000",
						 "000011000010000011111100",
						 "000011000010000000001000",
						 "000011000001111100010100",
						 "000011000001111000100000",
						 "000011000001110100101100",
						 "000011000001110000111000",
						 "000011000001101101000100",
						 "000011000001101001010000",
						 "000011000001100101011100",
						 "000011000001100001101000",
						 "000010111111110111110110",
						 "000010111111110100000010",
						 "000010111111110000001110",
						 "000010111111101100011010",
						 "000010111111101000100110",
						 "000010111111100100110010",
						 "000010111111100000111110",
						 "000010111111011101001010",
						 "000010111111011001010110",
						 "000010111111010101100010",
						 "000010111111010001101110",
						 "000010111111001101111010",
						 "000010111111001010000110",
						 "000010111111000110010010",
						 "000010111111000010011110",
						 "000010111110111110101010",
						 "000010111111110111110110",
						 "000010111111110100000010",
						 "000010111111110000001110",
						 "000010111111101100011010",
						 "000010111111101000100110",
						 "000010111111100100110010",
						 "000010111111100000111110",
						 "000010111111011101001010",
						 "000010111111011001010110",
						 "000010111111010101100010",
						 "000010111111010001101110",
						 "000010111111001101111010",
						 "000010111111001010000110",
						 "000010111111000110010010",
						 "000010111111000010011110",
						 "000010111110111110101010",
						 "000010111101010100111000",
						 "000010111101010001000100",
						 "000010111101001101010000",
						 "000010111101001001011100",
						 "000010111101000101101000",
						 "000010111101000001110100",
						 "000010111100111110000000",
						 "000010111100111010001100",
						 "000010111100110110011000",
						 "000010111100110010100100",
						 "000010111100101110110000",
						 "000010111100101010111100",
						 "000010111100100111001000",
						 "000010111100100011010100",
						 "000010111100011111100000",
						 "000010111100011011101100",
						 "000010111101010100111000",
						 "000010111101010001000100",
						 "000010111101001101010000",
						 "000010111101001001011100",
						 "000010111101000101101000",
						 "000010111101000001110100",
						 "000010111100111110000000",
						 "000010111100111010001100",
						 "000010111100110110011000",
						 "000010111100110010100100",
						 "000010111100101110110000",
						 "000010111100101010111100",
						 "000010111100100111001000",
						 "000010111100100011010100",
						 "000010111100011111100000",
						 "000010111100011011101100",
						 "000010111101010100111000",
						 "000010111101010001000100",
						 "000010111101001101010000",
						 "000010111101001001011100",
						 "000010111101000101101000",
						 "000010111101000001110100",
						 "000010111100111110000000",
						 "000010111100111010001100",
						 "000010111100110110011000",
						 "000010111100110010100100",
						 "000010111100101110110000",
						 "000010111100101010111100",
						 "000010111100100111001000",
						 "000010111100100011010100",
						 "000010111100011111100000",
						 "000010111100011011101100",
						 "000010111010110001111010",
						 "000010111010101110000110",
						 "000010111010101010010010",
						 "000010111010100110011110",
						 "000010111010100010101010",
						 "000010111010011110110110",
						 "000010111010011011000010",
						 "000010111010010111001110",
						 "000010111010010011011010",
						 "000010111010001111100110",
						 "000010111010001011110010",
						 "000010111010000111111110",
						 "000010111010000100001010",
						 "000010111010000000010110",
						 "000010111001111100100010",
						 "000010111001111000101110",
						 "000010111010110001111010",
						 "000010111010101110000110",
						 "000010111010101010010010",
						 "000010111010100110011110",
						 "000010111010100010101010",
						 "000010111010011110110110",
						 "000010111010011011000010",
						 "000010111010010111001110",
						 "000010111010010011011010",
						 "000010111010001111100110",
						 "000010111010001011110010",
						 "000010111010000111111110",
						 "000010111010000100001010",
						 "000010111010000000010110",
						 "000010111001111100100010",
						 "000010111001111000101110",
						 "000010111010110001111010",
						 "000010111010101110000110",
						 "000010111010101010010010",
						 "000010111010100110011110",
						 "000010111010100010101010",
						 "000010111010011110110110",
						 "000010111010011011000010",
						 "000010111010010111001110",
						 "000010111010010011011010",
						 "000010111010001111100110",
						 "000010111010001011110010",
						 "000010111010000111111110",
						 "000010111010000100001010",
						 "000010111010000000010110",
						 "000010111001111100100010",
						 "000010111001111000101110",
						 "000010111000001111001011",
						 "000010111000001011010110",
						 "000010111000000111100001",
						 "000010111000000011101100",
						 "000010110111111111110111",
						 "000010110111111100000010",
						 "000010110111111000001101",
						 "000010110111110100011000",
						 "000010110111110000100011",
						 "000010110111101100101110",
						 "000010110111101000111001",
						 "000010110111100101000100",
						 "000010110111100001001111",
						 "000010110111011101011010",
						 "000010110111011001100101",
						 "000010110111010101110000",
						 "000010111000001111001011",
						 "000010111000001011010110",
						 "000010111000000111100001",
						 "000010111000000011101100",
						 "000010110111111111110111",
						 "000010110111111100000010",
						 "000010110111111000001101",
						 "000010110111110100011000",
						 "000010110111110000100011",
						 "000010110111101100101110",
						 "000010110111101000111001",
						 "000010110111100101000100",
						 "000010110111100001001111",
						 "000010110111011101011010",
						 "000010110111011001100101",
						 "000010110111010101110000",
						 "000010110101101100001101",
						 "000010110101101000011000",
						 "000010110101100100100011",
						 "000010110101100000101110",
						 "000010110101011100111001",
						 "000010110101011001000100",
						 "000010110101010101001111",
						 "000010110101010001011010",
						 "000010110101001101100101",
						 "000010110101001001110000",
						 "000010110101000101111011",
						 "000010110101000010000110",
						 "000010110100111110010001",
						 "000010110100111010011100",
						 "000010110100110110100111",
						 "000010110100110010110010",
						 "000010110101101100001101",
						 "000010110101101000011000",
						 "000010110101100100100011",
						 "000010110101100000101110",
						 "000010110101011100111001",
						 "000010110101011001000100",
						 "000010110101010101001111",
						 "000010110101010001011010",
						 "000010110101001101100101",
						 "000010110101001001110000",
						 "000010110101000101111011",
						 "000010110101000010000110",
						 "000010110100111110010001",
						 "000010110100111010011100",
						 "000010110100110110100111",
						 "000010110100110010110010",
						 "000010110101101100001101",
						 "000010110101101000011000",
						 "000010110101100100100011",
						 "000010110101100000101110",
						 "000010110101011100111001",
						 "000010110101011001000100",
						 "000010110101010101001111",
						 "000010110101010001011010",
						 "000010110101001101100101",
						 "000010110101001001110000",
						 "000010110101000101111011",
						 "000010110101000010000110",
						 "000010110100111110010001",
						 "000010110100111010011100",
						 "000010110100110110100111",
						 "000010110100110010110010",
						 "000010110011001001001111",
						 "000010110011000101011010",
						 "000010110011000001100101",
						 "000010110010111101110000",
						 "000010110010111001111011",
						 "000010110010110110000110",
						 "000010110010110010010001",
						 "000010110010101110011100",
						 "000010110010101010100111",
						 "000010110010100110110010",
						 "000010110010100010111101",
						 "000010110010011111001000",
						 "000010110010011011010011",
						 "000010110010010111011110",
						 "000010110010010011101001",
						 "000010110010001111110100",
						 "000010110011001001001111",
						 "000010110011000101011010",
						 "000010110011000001100101",
						 "000010110010111101110000",
						 "000010110010111001111011",
						 "000010110010110110000110",
						 "000010110010110010010001",
						 "000010110010101110011100",
						 "000010110010101010100111",
						 "000010110010100110110010",
						 "000010110010100010111101",
						 "000010110010011111001000",
						 "000010110010011011010011",
						 "000010110010010111011110",
						 "000010110010010011101001",
						 "000010110010001111110100",
						 "000010110011001001001111",
						 "000010110011000101011010",
						 "000010110011000001100101",
						 "000010110010111101110000",
						 "000010110010111001111011",
						 "000010110010110110000110",
						 "000010110010110010010001",
						 "000010110010101110011100",
						 "000010110010101010100111",
						 "000010110010100110110010",
						 "000010110010100010111101",
						 "000010110010011111001000",
						 "000010110010011011010011",
						 "000010110010010111011110",
						 "000010110010010011101001",
						 "000010110010001111110100",
						 "000010110000100110010001",
						 "000010110000100010011100",
						 "000010110000011110100111",
						 "000010110000011010110010",
						 "000010110000010110111101",
						 "000010110000010011001000",
						 "000010110000001111010011",
						 "000010110000001011011110",
						 "000010110000000111101001",
						 "000010110000000011110100",
						 "000010101111111111111111",
						 "000010101111111100001010",
						 "000010101111111000010101",
						 "000010101111110100100000",
						 "000010101111110000101011",
						 "000010101111101100110110",
						 "000010110000100110010001",
						 "000010110000100010011100",
						 "000010110000011110100111",
						 "000010110000011010110010",
						 "000010110000010110111101",
						 "000010110000010011001000",
						 "000010110000001111010011",
						 "000010110000001011011110",
						 "000010110000000111101001",
						 "000010110000000011110100",
						 "000010101111111111111111",
						 "000010101111111100001010",
						 "000010101111111000010101",
						 "000010101111110100100000",
						 "000010101111110000101011",
						 "000010101111101100110110",
						 "000010101110000011100010",
						 "000010101101111111101100",
						 "000010101101111011110110",
						 "000010101101111000000000",
						 "000010101101110100001010",
						 "000010101101110000010100",
						 "000010101101101100011110",
						 "000010101101101000101000",
						 "000010101101100100110010",
						 "000010101101100000111100",
						 "000010101101011101000110",
						 "000010101101011001010000",
						 "000010101101010101011010",
						 "000010101101010001100100",
						 "000010101101001101101110",
						 "000010101101001001111000",
						 "000010101110000011100010",
						 "000010101101111111101100",
						 "000010101101111011110110",
						 "000010101101111000000000",
						 "000010101101110100001010",
						 "000010101101110000010100",
						 "000010101101101100011110",
						 "000010101101101000101000",
						 "000010101101100100110010",
						 "000010101101100000111100",
						 "000010101101011101000110",
						 "000010101101011001010000",
						 "000010101101010101011010",
						 "000010101101010001100100",
						 "000010101101001101101110",
						 "000010101101001001111000",
						 "000010101110000011100010",
						 "000010101101111111101100",
						 "000010101101111011110110",
						 "000010101101111000000000",
						 "000010101101110100001010",
						 "000010101101110000010100",
						 "000010101101101100011110",
						 "000010101101101000101000",
						 "000010101101100100110010",
						 "000010101101100000111100",
						 "000010101101011101000110",
						 "000010101101011001010000",
						 "000010101101010101011010",
						 "000010101101010001100100",
						 "000010101101001101101110",
						 "000010101101001001111000",
						 "000010101011100000100100",
						 "000010101011011100101110",
						 "000010101011011000111000",
						 "000010101011010101000010",
						 "000010101011010001001100",
						 "000010101011001101010110",
						 "000010101011001001100000",
						 "000010101011000101101010",
						 "000010101011000001110100",
						 "000010101010111101111110",
						 "000010101010111010001000",
						 "000010101010110110010010",
						 "000010101010110010011100",
						 "000010101010101110100110",
						 "000010101010101010110000",
						 "000010101010100110111010",
						 "000010101011100000100100",
						 "000010101011011100101110",
						 "000010101011011000111000",
						 "000010101011010101000010",
						 "000010101011010001001100",
						 "000010101011001101010110",
						 "000010101011001001100000",
						 "000010101011000101101010",
						 "000010101011000001110100",
						 "000010101010111101111110",
						 "000010101010111010001000",
						 "000010101010110110010010",
						 "000010101010110010011100",
						 "000010101010101110100110",
						 "000010101010101010110000",
						 "000010101010100110111010",
						 "000010101011100000100100",
						 "000010101011011100101110",
						 "000010101011011000111000",
						 "000010101011010101000010",
						 "000010101011010001001100",
						 "000010101011001101010110",
						 "000010101011001001100000",
						 "000010101011000101101010",
						 "000010101011000001110100",
						 "000010101010111101111110",
						 "000010101010111010001000",
						 "000010101010110110010010",
						 "000010101010110010011100",
						 "000010101010101110100110",
						 "000010101010101010110000",
						 "000010101010100110111010",
						 "000010101000111101100110",
						 "000010101000111001110000",
						 "000010101000110101111010",
						 "000010101000110010000100",
						 "000010101000101110001110",
						 "000010101000101010011000",
						 "000010101000100110100010",
						 "000010101000100010101100",
						 "000010101000011110110110",
						 "000010101000011011000000",
						 "000010101000010111001010",
						 "000010101000010011010100",
						 "000010101000001111011110",
						 "000010101000001011101000",
						 "000010101000000111110010",
						 "000010101000000011111100",
						 "000010101000111101100110",
						 "000010101000111001110000",
						 "000010101000110101111010",
						 "000010101000110010000100",
						 "000010101000101110001110",
						 "000010101000101010011000",
						 "000010101000100110100010",
						 "000010101000100010101100",
						 "000010101000011110110110",
						 "000010101000011011000000",
						 "000010101000010111001010",
						 "000010101000010011010100",
						 "000010101000001111011110",
						 "000010101000001011101000",
						 "000010101000000111110010",
						 "000010101000000011111100",
						 "000010100110011010101000",
						 "000010100110010110110010",
						 "000010100110010010111100",
						 "000010100110001111000110",
						 "000010100110001011010000",
						 "000010100110000111011010",
						 "000010100110000011100100",
						 "000010100101111111101110",
						 "000010100101111011111000",
						 "000010100101111000000010",
						 "000010100101110100001100",
						 "000010100101110000010110",
						 "000010100101101100100000",
						 "000010100101101000101010",
						 "000010100101100100110100",
						 "000010100101100000111110",
						 "000010100110011010110111",
						 "000010100110010111000000",
						 "000010100110010011001001",
						 "000010100110001111010010",
						 "000010100110001011011011",
						 "000010100110000111100100",
						 "000010100110000011101101",
						 "000010100101111111110110",
						 "000010100101111011111111",
						 "000010100101111000001000",
						 "000010100101110100010001",
						 "000010100101110000011010",
						 "000010100101101100100011",
						 "000010100101101000101100",
						 "000010100101100100110101",
						 "000010100101100000111110",
						 "000010100110011010110111",
						 "000010100110010111000000",
						 "000010100110010011001001",
						 "000010100110001111010010",
						 "000010100110001011011011",
						 "000010100110000111100100",
						 "000010100110000011101101",
						 "000010100101111111110110",
						 "000010100101111011111111",
						 "000010100101111000001000",
						 "000010100101110100010001",
						 "000010100101110000011010",
						 "000010100101101100100011",
						 "000010100101101000101100",
						 "000010100101100100110101",
						 "000010100101100000111110",
						 "000010100011110111111001",
						 "000010100011110100000010",
						 "000010100011110000001011",
						 "000010100011101100010100",
						 "000010100011101000011101",
						 "000010100011100100100110",
						 "000010100011100000101111",
						 "000010100011011100111000",
						 "000010100011011001000001",
						 "000010100011010101001010",
						 "000010100011010001010011",
						 "000010100011001101011100",
						 "000010100011001001100101",
						 "000010100011000101101110",
						 "000010100011000001110111",
						 "000010100010111110000000",
						 "000010100011110111111001",
						 "000010100011110100000010",
						 "000010100011110000001011",
						 "000010100011101100010100",
						 "000010100011101000011101",
						 "000010100011100100100110",
						 "000010100011100000101111",
						 "000010100011011100111000",
						 "000010100011011001000001",
						 "000010100011010101001010",
						 "000010100011010001010011",
						 "000010100011001101011100",
						 "000010100011001001100101",
						 "000010100011000101101110",
						 "000010100011000001110111",
						 "000010100010111110000000",
						 "000010100001010100111011",
						 "000010100001010001000100",
						 "000010100001001101001101",
						 "000010100001001001010110",
						 "000010100001000101011111",
						 "000010100001000001101000",
						 "000010100000111101110001",
						 "000010100000111001111010",
						 "000010100000110110000011",
						 "000010100000110010001100",
						 "000010100000101110010101",
						 "000010100000101010011110",
						 "000010100000100110100111",
						 "000010100000100010110000",
						 "000010100000011110111001",
						 "000010100000011011000010",
						 "000010100001010100111011",
						 "000010100001010001000100",
						 "000010100001001101001101",
						 "000010100001001001010110",
						 "000010100001000101011111",
						 "000010100001000001101000",
						 "000010100000111101110001",
						 "000010100000111001111010",
						 "000010100000110110000011",
						 "000010100000110010001100",
						 "000010100000101110010101",
						 "000010100000101010011110",
						 "000010100000100110100111",
						 "000010100000100010110000",
						 "000010100000011110111001",
						 "000010100000011011000010",
						 "000010100001010100111011",
						 "000010100001010001000100",
						 "000010100001001101001101",
						 "000010100001001001010110",
						 "000010100001000101011111",
						 "000010100001000001101000",
						 "000010100000111101110001",
						 "000010100000111001111010",
						 "000010100000110110000011",
						 "000010100000110010001100",
						 "000010100000101110010101",
						 "000010100000101010011110",
						 "000010100000100110100111",
						 "000010100000100010110000",
						 "000010100000011110111001",
						 "000010100000011011000010",
						 "000010011110110001111101",
						 "000010011110101110000110",
						 "000010011110101010001111",
						 "000010011110100110011000",
						 "000010011110100010100001",
						 "000010011110011110101010",
						 "000010011110011010110011",
						 "000010011110010110111100",
						 "000010011110010011000101",
						 "000010011110001111001110",
						 "000010011110001011010111",
						 "000010011110000111100000",
						 "000010011110000011101001",
						 "000010011101111111110010",
						 "000010011101111011111011",
						 "000010011101111000000100",
						 "000010011110110001111101",
						 "000010011110101110000110",
						 "000010011110101010001111",
						 "000010011110100110011000",
						 "000010011110100010100001",
						 "000010011110011110101010",
						 "000010011110011010110011",
						 "000010011110010110111100",
						 "000010011110010011000101",
						 "000010011110001111001110",
						 "000010011110001011010111",
						 "000010011110000111100000",
						 "000010011110000011101001",
						 "000010011101111111110010",
						 "000010011101111011111011",
						 "000010011101111000000100",
						 "000010011110110001111101",
						 "000010011110101110000110",
						 "000010011110101010001111",
						 "000010011110100110011000",
						 "000010011110100010100001",
						 "000010011110011110101010",
						 "000010011110011010110011",
						 "000010011110010110111100",
						 "000010011110010011000101",
						 "000010011110001111001110",
						 "000010011110001011010111",
						 "000010011110000111100000",
						 "000010011110000011101001",
						 "000010011101111111110010",
						 "000010011101111011111011",
						 "000010011101111000000100",
						 "000010011100001110111111",
						 "000010011100001011001000",
						 "000010011100000111010001",
						 "000010011100000011011010",
						 "000010011011111111100011",
						 "000010011011111011101100",
						 "000010011011110111110101",
						 "000010011011110011111110",
						 "000010011011110000000111",
						 "000010011011101100010000",
						 "000010011011101000011001",
						 "000010011011100100100010",
						 "000010011011100000101011",
						 "000010011011011100110100",
						 "000010011011011000111101",
						 "000010011011010101000110",
						 "000010011100001111001110",
						 "000010011100001011010110",
						 "000010011100000111011110",
						 "000010011100000011100110",
						 "000010011011111111101110",
						 "000010011011111011110110",
						 "000010011011110111111110",
						 "000010011011110100000110",
						 "000010011011110000001110",
						 "000010011011101100010110",
						 "000010011011101000011110",
						 "000010011011100100100110",
						 "000010011011100000101110",
						 "000010011011011100110110",
						 "000010011011011000111110",
						 "000010011011010101000110",
						 "000010011001101100010000",
						 "000010011001101000011000",
						 "000010011001100100100000",
						 "000010011001100000101000",
						 "000010011001011100110000",
						 "000010011001011000111000",
						 "000010011001010101000000",
						 "000010011001010001001000",
						 "000010011001001101010000",
						 "000010011001001001011000",
						 "000010011001000101100000",
						 "000010011001000001101000",
						 "000010011000111101110000",
						 "000010011000111001111000",
						 "000010011000110110000000",
						 "000010011000110010001000",
						 "000010011001101100010000",
						 "000010011001101000011000",
						 "000010011001100100100000",
						 "000010011001100000101000",
						 "000010011001011100110000",
						 "000010011001011000111000",
						 "000010011001010101000000",
						 "000010011001010001001000",
						 "000010011001001101010000",
						 "000010011001001001011000",
						 "000010011001000101100000",
						 "000010011001000001101000",
						 "000010011000111101110000",
						 "000010011000111001111000",
						 "000010011000110110000000",
						 "000010011000110010001000",
						 "000010011001101100010000",
						 "000010011001101000011000",
						 "000010011001100100100000",
						 "000010011001100000101000",
						 "000010011001011100110000",
						 "000010011001011000111000",
						 "000010011001010101000000",
						 "000010011001010001001000",
						 "000010011001001101010000",
						 "000010011001001001011000",
						 "000010011001000101100000",
						 "000010011001000001101000",
						 "000010011000111101110000",
						 "000010011000111001111000",
						 "000010011000110110000000",
						 "000010011000110010001000",
						 "000010010111001001010010",
						 "000010010111000101011010",
						 "000010010111000001100010",
						 "000010010110111101101010",
						 "000010010110111001110010",
						 "000010010110110101111010",
						 "000010010110110010000010",
						 "000010010110101110001010",
						 "000010010110101010010010",
						 "000010010110100110011010",
						 "000010010110100010100010",
						 "000010010110011110101010",
						 "000010010110011010110010",
						 "000010010110010110111010",
						 "000010010110010011000010",
						 "000010010110001111001010",
						 "000010010111001001010010",
						 "000010010111000101011010",
						 "000010010111000001100010",
						 "000010010110111101101010",
						 "000010010110111001110010",
						 "000010010110110101111010",
						 "000010010110110010000010",
						 "000010010110101110001010",
						 "000010010110101010010010",
						 "000010010110100110011010",
						 "000010010110100010100010",
						 "000010010110011110101010",
						 "000010010110011010110010",
						 "000010010110010110111010",
						 "000010010110010011000010",
						 "000010010110001111001010",
						 "000010010111001001010010",
						 "000010010111000101011010",
						 "000010010111000001100010",
						 "000010010110111101101010",
						 "000010010110111001110010",
						 "000010010110110101111010",
						 "000010010110110010000010",
						 "000010010110101110001010",
						 "000010010110101010010010",
						 "000010010110100110011010",
						 "000010010110100010100010",
						 "000010010110011110101010",
						 "000010010110011010110010",
						 "000010010110010110111010",
						 "000010010110010011000010",
						 "000010010110001111001010",
						 "000010010100100110010100",
						 "000010010100100010011100",
						 "000010010100011110100100",
						 "000010010100011010101100",
						 "000010010100010110110100",
						 "000010010100010010111100",
						 "000010010100001111000100",
						 "000010010100001011001100",
						 "000010010100000111010100",
						 "000010010100000011011100",
						 "000010010011111111100100",
						 "000010010011111011101100",
						 "000010010011110111110100",
						 "000010010011110011111100",
						 "000010010011110000000100",
						 "000010010011101100001100",
						 "000010010100100110010100",
						 "000010010100100010011100",
						 "000010010100011110100100",
						 "000010010100011010101100",
						 "000010010100010110110100",
						 "000010010100010010111100",
						 "000010010100001111000100",
						 "000010010100001011001100",
						 "000010010100000111010100",
						 "000010010100000011011100",
						 "000010010011111111100100",
						 "000010010011111011101100",
						 "000010010011110111110100",
						 "000010010011110011111100",
						 "000010010011110000000100",
						 "000010010011101100001100",
						 "000010010010000011010110",
						 "000010010001111111011110",
						 "000010010001111011100110",
						 "000010010001110111101110",
						 "000010010001110011110110",
						 "000010010001101111111110",
						 "000010010001101100000110",
						 "000010010001101000001110",
						 "000010010001100100010110",
						 "000010010001100000011110",
						 "000010010001011100100110",
						 "000010010001011000101110",
						 "000010010001010100110110",
						 "000010010001010000111110",
						 "000010010001001101000110",
						 "000010010001001001001110",
						 "000010010010000011100101",
						 "000010010001111111101100",
						 "000010010001111011110011",
						 "000010010001110111111010",
						 "000010010001110100000001",
						 "000010010001110000001000",
						 "000010010001101100001111",
						 "000010010001101000010110",
						 "000010010001100100011101",
						 "000010010001100000100100",
						 "000010010001011100101011",
						 "000010010001011000110010",
						 "000010010001010100111001",
						 "000010010001010001000000",
						 "000010010001001101000111",
						 "000010010001001001001110",
						 "000010010010000011100101",
						 "000010010001111111101100",
						 "000010010001111011110011",
						 "000010010001110111111010",
						 "000010010001110100000001",
						 "000010010001110000001000",
						 "000010010001101100001111",
						 "000010010001101000010110",
						 "000010010001100100011101",
						 "000010010001100000100100",
						 "000010010001011100101011",
						 "000010010001011000110010",
						 "000010010001010100111001",
						 "000010010001010001000000",
						 "000010010001001101000111",
						 "000010010001001001001110",
						 "000010001111100000100111",
						 "000010001111011100101110",
						 "000010001111011000110101",
						 "000010001111010100111100",
						 "000010001111010001000011",
						 "000010001111001101001010",
						 "000010001111001001010001",
						 "000010001111000101011000",
						 "000010001111000001011111",
						 "000010001110111101100110",
						 "000010001110111001101101",
						 "000010001110110101110100",
						 "000010001110110001111011",
						 "000010001110101110000010",
						 "000010001110101010001001",
						 "000010001110100110010000",
						 "000010001111100000100111",
						 "000010001111011100101110",
						 "000010001111011000110101",
						 "000010001111010100111100",
						 "000010001111010001000011",
						 "000010001111001101001010",
						 "000010001111001001010001",
						 "000010001111000101011000",
						 "000010001111000001011111",
						 "000010001110111101100110",
						 "000010001110111001101101",
						 "000010001110110101110100",
						 "000010001110110001111011",
						 "000010001110101110000010",
						 "000010001110101010001001",
						 "000010001110100110010000",
						 "000010001100111101101001",
						 "000010001100111001110000",
						 "000010001100110101110111",
						 "000010001100110001111110",
						 "000010001100101110000101",
						 "000010001100101010001100",
						 "000010001100100110010011",
						 "000010001100100010011010",
						 "000010001100011110100001",
						 "000010001100011010101000",
						 "000010001100010110101111",
						 "000010001100010010110110",
						 "000010001100001110111101",
						 "000010001100001011000100",
						 "000010001100000111001011",
						 "000010001100000011010010",
						 "000010001100111101101001",
						 "000010001100111001110000",
						 "000010001100110101110111",
						 "000010001100110001111110",
						 "000010001100101110000101",
						 "000010001100101010001100",
						 "000010001100100110010011",
						 "000010001100100010011010",
						 "000010001100011110100001",
						 "000010001100011010101000",
						 "000010001100010110101111",
						 "000010001100010010110110",
						 "000010001100001110111101",
						 "000010001100001011000100",
						 "000010001100000111001011",
						 "000010001100000011010010",
						 "000010001100111101101001",
						 "000010001100111001110000",
						 "000010001100110101110111",
						 "000010001100110001111110",
						 "000010001100101110000101",
						 "000010001100101010001100",
						 "000010001100100110010011",
						 "000010001100100010011010",
						 "000010001100011110100001",
						 "000010001100011010101000",
						 "000010001100010110101111",
						 "000010001100010010110110",
						 "000010001100001110111101",
						 "000010001100001011000100",
						 "000010001100000111001011",
						 "000010001100000011010010",
						 "000010001010011010101011",
						 "000010001010010110110010",
						 "000010001010010010111001",
						 "000010001010001111000000",
						 "000010001010001011000111",
						 "000010001010000111001110",
						 "000010001010000011010101",
						 "000010001001111111011100",
						 "000010001001111011100011",
						 "000010001001110111101010",
						 "000010001001110011110001",
						 "000010001001101111111000",
						 "000010001001101011111111",
						 "000010001001101000000110",
						 "000010001001100100001101",
						 "000010001001100000010100",
						 "000010001010011010101011",
						 "000010001010010110110010",
						 "000010001010010010111001",
						 "000010001010001111000000",
						 "000010001010001011000111",
						 "000010001010000111001110",
						 "000010001010000011010101",
						 "000010001001111111011100",
						 "000010001001111011100011",
						 "000010001001110111101010",
						 "000010001001110011110001",
						 "000010001001101111111000",
						 "000010001001101011111111",
						 "000010001001101000000110",
						 "000010001001100100001101",
						 "000010001001100000010100",
						 "000010001010011010101011",
						 "000010001010010110110010",
						 "000010001010010010111001",
						 "000010001010001111000000",
						 "000010001010001011000111",
						 "000010001010000111001110",
						 "000010001010000011010101",
						 "000010001001111111011100",
						 "000010001001111011100011",
						 "000010001001110111101010",
						 "000010001001110011110001",
						 "000010001001101111111000",
						 "000010001001101011111111",
						 "000010001001101000000110",
						 "000010001001100100001101",
						 "000010001001100000010100",
						 "000010000111110111101101",
						 "000010000111110011110100",
						 "000010000111101111111011",
						 "000010000111101100000010",
						 "000010000111101000001001",
						 "000010000111100100010000",
						 "000010000111100000010111",
						 "000010000111011100011110",
						 "000010000111011000100101",
						 "000010000111010100101100",
						 "000010000111010000110011",
						 "000010000111001100111010",
						 "000010000111001001000001",
						 "000010000111000101001000",
						 "000010000111000001001111",
						 "000010000110111101010110",
						 "000010000111110111101101",
						 "000010000111110011110100",
						 "000010000111101111111011",
						 "000010000111101100000010",
						 "000010000111101000001001",
						 "000010000111100100010000",
						 "000010000111100000010111",
						 "000010000111011100011110",
						 "000010000111011000100101",
						 "000010000111010100101100",
						 "000010000111010000110011",
						 "000010000111001100111010",
						 "000010000111001001000001",
						 "000010000111000101001000",
						 "000010000111000001001111",
						 "000010000110111101010110",
						 "000010000101010100111110",
						 "000010000101010001000100",
						 "000010000101001101001010",
						 "000010000101001001010000",
						 "000010000101000101010110",
						 "000010000101000001011100",
						 "000010000100111101100010",
						 "000010000100111001101000",
						 "000010000100110101101110",
						 "000010000100110001110100",
						 "000010000100101101111010",
						 "000010000100101010000000",
						 "000010000100100110000110",
						 "000010000100100010001100",
						 "000010000100011110010010",
						 "000010000100011010011000",
						 "000010000101010100111110",
						 "000010000101010001000100",
						 "000010000101001101001010",
						 "000010000101001001010000",
						 "000010000101000101010110",
						 "000010000101000001011100",
						 "000010000100111101100010",
						 "000010000100111001101000",
						 "000010000100110101101110",
						 "000010000100110001110100",
						 "000010000100101101111010",
						 "000010000100101010000000",
						 "000010000100100110000110",
						 "000010000100100010001100",
						 "000010000100011110010010",
						 "000010000100011010011000",
						 "000010000101010100111110",
						 "000010000101010001000100",
						 "000010000101001101001010",
						 "000010000101001001010000",
						 "000010000101000101010110",
						 "000010000101000001011100",
						 "000010000100111101100010",
						 "000010000100111001101000",
						 "000010000100110101101110",
						 "000010000100110001110100",
						 "000010000100101101111010",
						 "000010000100101010000000",
						 "000010000100100110000110",
						 "000010000100100010001100",
						 "000010000100011110010010",
						 "000010000100011010011000",
						 "000010000010110010000000",
						 "000010000010101110000110",
						 "000010000010101010001100",
						 "000010000010100110010010",
						 "000010000010100010011000",
						 "000010000010011110011110",
						 "000010000010011010100100",
						 "000010000010010110101010",
						 "000010000010010010110000",
						 "000010000010001110110110",
						 "000010000010001010111100",
						 "000010000010000111000010",
						 "000010000010000011001000",
						 "000010000001111111001110",
						 "000010000001111011010100",
						 "000010000001110111011010",
						 "000010000010110010000000",
						 "000010000010101110000110",
						 "000010000010101010001100",
						 "000010000010100110010010",
						 "000010000010100010011000",
						 "000010000010011110011110",
						 "000010000010011010100100",
						 "000010000010010110101010",
						 "000010000010010010110000",
						 "000010000010001110110110",
						 "000010000010001010111100",
						 "000010000010000111000010",
						 "000010000010000011001000",
						 "000010000001111111001110",
						 "000010000001111011010100",
						 "000010000001110111011010",
						 "000010000010110010000000",
						 "000010000010101110000110",
						 "000010000010101010001100",
						 "000010000010100110010010",
						 "000010000010100010011000",
						 "000010000010011110011110",
						 "000010000010011010100100",
						 "000010000010010110101010",
						 "000010000010010010110000",
						 "000010000010001110110110",
						 "000010000010001010111100",
						 "000010000010000111000010",
						 "000010000010000011001000",
						 "000010000001111111001110",
						 "000010000001111011010100",
						 "000010000001110111011010",
						 "000010000000001111000010",
						 "000010000000001011001000",
						 "000010000000000111001110",
						 "000010000000000011010100",
						 "000001111111111111011010",
						 "000001111111111011100000",
						 "000001111111110111100110",
						 "000001111111110011101100",
						 "000001111111101111110010",
						 "000001111111101011111000",
						 "000001111111100111111110",
						 "000001111111100100000100",
						 "000001111111100000001010",
						 "000001111111011100010000",
						 "000001111111011000010110",
						 "000001111111010100011100",
						 "000010000000001111000010",
						 "000010000000001011001000",
						 "000010000000000111001110",
						 "000010000000000011010100",
						 "000001111111111111011010",
						 "000001111111111011100000",
						 "000001111111110111100110",
						 "000001111111110011101100",
						 "000001111111101111110010",
						 "000001111111101011111000",
						 "000001111111100111111110",
						 "000001111111100100000100",
						 "000001111111100000001010",
						 "000001111111011100010000",
						 "000001111111011000010110",
						 "000001111111010100011100",
						 "000001111101101100000100",
						 "000001111101101000001010",
						 "000001111101100100010000",
						 "000001111101100000010110",
						 "000001111101011100011100",
						 "000001111101011000100010",
						 "000001111101010100101000",
						 "000001111101010000101110",
						 "000001111101001100110100",
						 "000001111101001000111010",
						 "000001111101000101000000",
						 "000001111101000001000110",
						 "000001111100111101001100",
						 "000001111100111001010010",
						 "000001111100110101011000",
						 "000001111100110001011110",
						 "000001111101101100000100",
						 "000001111101101000001010",
						 "000001111101100100010000",
						 "000001111101100000010110",
						 "000001111101011100011100",
						 "000001111101011000100010",
						 "000001111101010100101000",
						 "000001111101010000101110",
						 "000001111101001100110100",
						 "000001111101001000111010",
						 "000001111101000101000000",
						 "000001111101000001000110",
						 "000001111100111101001100",
						 "000001111100111001010010",
						 "000001111100110101011000",
						 "000001111100110001011110",
						 "000001111101101100000100",
						 "000001111101101000001010",
						 "000001111101100100010000",
						 "000001111101100000010110",
						 "000001111101011100011100",
						 "000001111101011000100010",
						 "000001111101010100101000",
						 "000001111101010000101110",
						 "000001111101001100110100",
						 "000001111101001000111010",
						 "000001111101000101000000",
						 "000001111101000001000110",
						 "000001111100111101001100",
						 "000001111100111001010010",
						 "000001111100110101011000",
						 "000001111100110001011110",
						 "000001111011001001000110",
						 "000001111011000101001100",
						 "000001111011000001010010",
						 "000001111010111101011000",
						 "000001111010111001011110",
						 "000001111010110101100100",
						 "000001111010110001101010",
						 "000001111010101101110000",
						 "000001111010101001110110",
						 "000001111010100101111100",
						 "000001111010100010000010",
						 "000001111010011110001000",
						 "000001111010011010001110",
						 "000001111010010110010100",
						 "000001111010010010011010",
						 "000001111010001110100000",
						 "000001111011001001000110",
						 "000001111011000101001100",
						 "000001111011000001010010",
						 "000001111010111101011000",
						 "000001111010111001011110",
						 "000001111010110101100100",
						 "000001111010110001101010",
						 "000001111010101101110000",
						 "000001111010101001110110",
						 "000001111010100101111100",
						 "000001111010100010000010",
						 "000001111010011110001000",
						 "000001111010011010001110",
						 "000001111010010110010100",
						 "000001111010010010011010",
						 "000001111010001110100000",
						 "000001111000100110010111",
						 "000001111000100010011100",
						 "000001111000011110100001",
						 "000001111000011010100110",
						 "000001111000010110101011",
						 "000001111000010010110000",
						 "000001111000001110110101",
						 "000001111000001010111010",
						 "000001111000000110111111",
						 "000001111000000011000100",
						 "000001110111111111001001",
						 "000001110111111011001110",
						 "000001110111110111010011",
						 "000001110111110011011000",
						 "000001110111101111011101",
						 "000001110111101011100010",
						 "000001111000100110010111",
						 "000001111000100010011100",
						 "000001111000011110100001",
						 "000001111000011010100110",
						 "000001111000010110101011",
						 "000001111000010010110000",
						 "000001111000001110110101",
						 "000001111000001010111010",
						 "000001111000000110111111",
						 "000001111000000011000100",
						 "000001110111111111001001",
						 "000001110111111011001110",
						 "000001110111110111010011",
						 "000001110111110011011000",
						 "000001110111101111011101",
						 "000001110111101011100010",
						 "000001111000100110010111",
						 "000001111000100010011100",
						 "000001111000011110100001",
						 "000001111000011010100110",
						 "000001111000010110101011",
						 "000001111000010010110000",
						 "000001111000001110110101",
						 "000001111000001010111010",
						 "000001111000000110111111",
						 "000001111000000011000100",
						 "000001110111111111001001",
						 "000001110111111011001110",
						 "000001110111110111010011",
						 "000001110111110011011000",
						 "000001110111101111011101",
						 "000001110111101011100010",
						 "000001110110000011011001",
						 "000001110101111111011110",
						 "000001110101111011100011",
						 "000001110101110111101000",
						 "000001110101110011101101",
						 "000001110101101111110010",
						 "000001110101101011110111",
						 "000001110101100111111100",
						 "000001110101100100000001",
						 "000001110101100000000110",
						 "000001110101011100001011",
						 "000001110101011000010000",
						 "000001110101010100010101",
						 "000001110101010000011010",
						 "000001110101001100011111",
						 "000001110101001000100100",
						 "000001110110000011011001",
						 "000001110101111111011110",
						 "000001110101111011100011",
						 "000001110101110111101000",
						 "000001110101110011101101",
						 "000001110101101111110010",
						 "000001110101101011110111",
						 "000001110101100111111100",
						 "000001110101100100000001",
						 "000001110101100000000110",
						 "000001110101011100001011",
						 "000001110101011000010000",
						 "000001110101010100010101",
						 "000001110101010000011010",
						 "000001110101001100011111",
						 "000001110101001000100100",
						 "000001110110000011011001",
						 "000001110101111111011110",
						 "000001110101111011100011",
						 "000001110101110111101000",
						 "000001110101110011101101",
						 "000001110101101111110010",
						 "000001110101101011110111",
						 "000001110101100111111100",
						 "000001110101100100000001",
						 "000001110101100000000110",
						 "000001110101011100001011",
						 "000001110101011000010000",
						 "000001110101010100010101",
						 "000001110101010000011010",
						 "000001110101001100011111",
						 "000001110101001000100100",
						 "000001110011100000011011",
						 "000001110011011100100000",
						 "000001110011011000100101",
						 "000001110011010100101010",
						 "000001110011010000101111",
						 "000001110011001100110100",
						 "000001110011001000111001",
						 "000001110011000100111110",
						 "000001110011000001000011",
						 "000001110010111101001000",
						 "000001110010111001001101",
						 "000001110010110101010010",
						 "000001110010110001010111",
						 "000001110010101101011100",
						 "000001110010101001100001",
						 "000001110010100101100110",
						 "000001110011100000011011",
						 "000001110011011100100000",
						 "000001110011011000100101",
						 "000001110011010100101010",
						 "000001110011010000101111",
						 "000001110011001100110100",
						 "000001110011001000111001",
						 "000001110011000100111110",
						 "000001110011000001000011",
						 "000001110010111101001000",
						 "000001110010111001001101",
						 "000001110010110101010010",
						 "000001110010110001010111",
						 "000001110010101101011100",
						 "000001110010101001100001",
						 "000001110010100101100110",
						 "000001110000111101011101",
						 "000001110000111001100010",
						 "000001110000110101100111",
						 "000001110000110001101100",
						 "000001110000101101110001",
						 "000001110000101001110110",
						 "000001110000100101111011",
						 "000001110000100010000000",
						 "000001110000011110000101",
						 "000001110000011010001010",
						 "000001110000010110001111",
						 "000001110000010010010100",
						 "000001110000001110011001",
						 "000001110000001010011110",
						 "000001110000000110100011",
						 "000001110000000010101000",
						 "000001110000111101011101",
						 "000001110000111001100010",
						 "000001110000110101100111",
						 "000001110000110001101100",
						 "000001110000101101110001",
						 "000001110000101001110110",
						 "000001110000100101111011",
						 "000001110000100010000000",
						 "000001110000011110000101",
						 "000001110000011010001010",
						 "000001110000010110001111",
						 "000001110000010010010100",
						 "000001110000001110011001",
						 "000001110000001010011110",
						 "000001110000000110100011",
						 "000001110000000010101000",
						 "000001110000111101011101",
						 "000001110000111001100010",
						 "000001110000110101100111",
						 "000001110000110001101100",
						 "000001110000101101110001",
						 "000001110000101001110110",
						 "000001110000100101111011",
						 "000001110000100010000000",
						 "000001110000011110000101",
						 "000001110000011010001010",
						 "000001110000010110001111",
						 "000001110000010010010100",
						 "000001110000001110011001",
						 "000001110000001010011110",
						 "000001110000000110100011",
						 "000001110000000010101000",
						 "000001101110011010011111",
						 "000001101110010110100100",
						 "000001101110010010101001",
						 "000001101110001110101110",
						 "000001101110001010110011",
						 "000001101110000110111000",
						 "000001101110000010111101",
						 "000001101101111111000010",
						 "000001101101111011000111",
						 "000001101101110111001100",
						 "000001101101110011010001",
						 "000001101101101111010110",
						 "000001101101101011011011",
						 "000001101101100111100000",
						 "000001101101100011100101",
						 "000001101101011111101010",
						 "000001101110011010011111",
						 "000001101110010110100100",
						 "000001101110010010101001",
						 "000001101110001110101110",
						 "000001101110001010110011",
						 "000001101110000110111000",
						 "000001101110000010111101",
						 "000001101101111111000010",
						 "000001101101111011000111",
						 "000001101101110111001100",
						 "000001101101110011010001",
						 "000001101101101111010110",
						 "000001101101101011011011",
						 "000001101101100111100000",
						 "000001101101100011100101",
						 "000001101101011111101010",
						 "000001101011110111100001",
						 "000001101011110011100110",
						 "000001101011101111101011",
						 "000001101011101011110000",
						 "000001101011100111110101",
						 "000001101011100011111010",
						 "000001101011011111111111",
						 "000001101011011100000100",
						 "000001101011011000001001",
						 "000001101011010100001110",
						 "000001101011010000010011",
						 "000001101011001100011000",
						 "000001101011001000011101",
						 "000001101011000100100010",
						 "000001101011000000100111",
						 "000001101010111100101100",
						 "000001101011110111100001",
						 "000001101011110011100110",
						 "000001101011101111101011",
						 "000001101011101011110000",
						 "000001101011100111110101",
						 "000001101011100011111010",
						 "000001101011011111111111",
						 "000001101011011100000100",
						 "000001101011011000001001",
						 "000001101011010100001110",
						 "000001101011010000010011",
						 "000001101011001100011000",
						 "000001101011001000011101",
						 "000001101011000100100010",
						 "000001101011000000100111",
						 "000001101010111100101100",
						 "000001101011110111110000",
						 "000001101011110011110100",
						 "000001101011101111111000",
						 "000001101011101011111100",
						 "000001101011101000000000",
						 "000001101011100100000100",
						 "000001101011100000001000",
						 "000001101011011100001100",
						 "000001101011011000010000",
						 "000001101011010100010100",
						 "000001101011010000011000",
						 "000001101011001100011100",
						 "000001101011001000100000",
						 "000001101011000100100100",
						 "000001101011000000101000",
						 "000001101010111100101100",
						 "000001101001010100110010",
						 "000001101001010000110110",
						 "000001101001001100111010",
						 "000001101001001000111110",
						 "000001101001000101000010",
						 "000001101001000001000110",
						 "000001101000111101001010",
						 "000001101000111001001110",
						 "000001101000110101010010",
						 "000001101000110001010110",
						 "000001101000101101011010",
						 "000001101000101001011110",
						 "000001101000100101100010",
						 "000001101000100001100110",
						 "000001101000011101101010",
						 "000001101000011001101110",
						 "000001101001010100110010",
						 "000001101001010000110110",
						 "000001101001001100111010",
						 "000001101001001000111110",
						 "000001101001000101000010",
						 "000001101001000001000110",
						 "000001101000111101001010",
						 "000001101000111001001110",
						 "000001101000110101010010",
						 "000001101000110001010110",
						 "000001101000101101011010",
						 "000001101000101001011110",
						 "000001101000100101100010",
						 "000001101000100001100110",
						 "000001101000011101101010",
						 "000001101000011001101110",
						 "000001101001010100110010",
						 "000001101001010000110110",
						 "000001101001001100111010",
						 "000001101001001000111110",
						 "000001101001000101000010",
						 "000001101001000001000110",
						 "000001101000111101001010",
						 "000001101000111001001110",
						 "000001101000110101010010",
						 "000001101000110001010110",
						 "000001101000101101011010",
						 "000001101000101001011110",
						 "000001101000100101100010",
						 "000001101000100001100110",
						 "000001101000011101101010",
						 "000001101000011001101110",
						 "000001100110110001110100",
						 "000001100110101101111000",
						 "000001100110101001111100",
						 "000001100110100110000000",
						 "000001100110100010000100",
						 "000001100110011110001000",
						 "000001100110011010001100",
						 "000001100110010110010000",
						 "000001100110010010010100",
						 "000001100110001110011000",
						 "000001100110001010011100",
						 "000001100110000110100000",
						 "000001100110000010100100",
						 "000001100101111110101000",
						 "000001100101111010101100",
						 "000001100101110110110000",
						 "000001100110110001110100",
						 "000001100110101101111000",
						 "000001100110101001111100",
						 "000001100110100110000000",
						 "000001100110100010000100",
						 "000001100110011110001000",
						 "000001100110011010001100",
						 "000001100110010110010000",
						 "000001100110010010010100",
						 "000001100110001110011000",
						 "000001100110001010011100",
						 "000001100110000110100000",
						 "000001100110000010100100",
						 "000001100101111110101000",
						 "000001100101111010101100",
						 "000001100101110110110000",
						 "000001100100001110110110",
						 "000001100100001010111010",
						 "000001100100000110111110",
						 "000001100100000011000010",
						 "000001100011111111000110",
						 "000001100011111011001010",
						 "000001100011110111001110",
						 "000001100011110011010010",
						 "000001100011101111010110",
						 "000001100011101011011010",
						 "000001100011100111011110",
						 "000001100011100011100010",
						 "000001100011011111100110",
						 "000001100011011011101010",
						 "000001100011010111101110",
						 "000001100011010011110010",
						 "000001100100001110110110",
						 "000001100100001010111010",
						 "000001100100000110111110",
						 "000001100100000011000010",
						 "000001100011111111000110",
						 "000001100011111011001010",
						 "000001100011110111001110",
						 "000001100011110011010010",
						 "000001100011101111010110",
						 "000001100011101011011010",
						 "000001100011100111011110",
						 "000001100011100011100010",
						 "000001100011011111100110",
						 "000001100011011011101010",
						 "000001100011010111101110",
						 "000001100011010011110010",
						 "000001100100001110110110",
						 "000001100100001010111010",
						 "000001100100000110111110",
						 "000001100100000011000010",
						 "000001100011111111000110",
						 "000001100011111011001010",
						 "000001100011110111001110",
						 "000001100011110011010010",
						 "000001100011101111010110",
						 "000001100011101011011010",
						 "000001100011100111011110",
						 "000001100011100011100010",
						 "000001100011011111100110",
						 "000001100011011011101010",
						 "000001100011010111101110",
						 "000001100011010011110010",
						 "000001100001101011111000",
						 "000001100001100111111100",
						 "000001100001100100000000",
						 "000001100001100000000100",
						 "000001100001011100001000",
						 "000001100001011000001100",
						 "000001100001010100010000",
						 "000001100001010000010100",
						 "000001100001001100011000",
						 "000001100001001000011100",
						 "000001100001000100100000",
						 "000001100001000000100100",
						 "000001100000111100101000",
						 "000001100000111000101100",
						 "000001100000110100110000",
						 "000001100000110000110100",
						 "000001100001101011111000",
						 "000001100001100111111100",
						 "000001100001100100000000",
						 "000001100001100000000100",
						 "000001100001011100001000",
						 "000001100001011000001100",
						 "000001100001010100010000",
						 "000001100001010000010100",
						 "000001100001001100011000",
						 "000001100001001000011100",
						 "000001100001000100100000",
						 "000001100001000000100100",
						 "000001100000111100101000",
						 "000001100000111000101100",
						 "000001100000110100110000",
						 "000001100000110000110100",
						 "000001011111001000111010",
						 "000001011111000100111110",
						 "000001011111000001000010",
						 "000001011110111101000110",
						 "000001011110111001001010",
						 "000001011110110101001110",
						 "000001011110110001010010",
						 "000001011110101101010110",
						 "000001011110101001011010",
						 "000001011110100101011110",
						 "000001011110100001100010",
						 "000001011110011101100110",
						 "000001011110011001101010",
						 "000001011110010101101110",
						 "000001011110010001110010",
						 "000001011110001101110110",
						 "000001011111001000111010",
						 "000001011111000100111110",
						 "000001011111000001000010",
						 "000001011110111101000110",
						 "000001011110111001001010",
						 "000001011110110101001110",
						 "000001011110110001010010",
						 "000001011110101101010110",
						 "000001011110101001011010",
						 "000001011110100101011110",
						 "000001011110100001100010",
						 "000001011110011101100110",
						 "000001011110011001101010",
						 "000001011110010101101110",
						 "000001011110010001110010",
						 "000001011110001101110110",
						 "000001011111001000111010",
						 "000001011111000100111110",
						 "000001011111000001000010",
						 "000001011110111101000110",
						 "000001011110111001001010",
						 "000001011110110101001110",
						 "000001011110110001010010",
						 "000001011110101101010110",
						 "000001011110101001011010",
						 "000001011110100101011110",
						 "000001011110100001100010",
						 "000001011110011101100110",
						 "000001011110011001101010",
						 "000001011110010101101110",
						 "000001011110010001110010",
						 "000001011110001101110110",
						 "000001011100100101111100",
						 "000001011100100010000000",
						 "000001011100011110000100",
						 "000001011100011010001000",
						 "000001011100010110001100",
						 "000001011100010010010000",
						 "000001011100001110010100",
						 "000001011100001010011000",
						 "000001011100000110011100",
						 "000001011100000010100000",
						 "000001011011111110100100",
						 "000001011011111010101000",
						 "000001011011110110101100",
						 "000001011011110010110000",
						 "000001011011101110110100",
						 "000001011011101010111000",
						 "000001011100100101111100",
						 "000001011100100010000000",
						 "000001011100011110000100",
						 "000001011100011010001000",
						 "000001011100010110001100",
						 "000001011100010010010000",
						 "000001011100001110010100",
						 "000001011100001010011000",
						 "000001011100000110011100",
						 "000001011100000010100000",
						 "000001011011111110100100",
						 "000001011011111010101000",
						 "000001011011110110101100",
						 "000001011011110010110000",
						 "000001011011101110110100",
						 "000001011011101010111000",
						 "000001011010000010111110",
						 "000001011001111111000010",
						 "000001011001111011000110",
						 "000001011001110111001010",
						 "000001011001110011001110",
						 "000001011001101111010010",
						 "000001011001101011010110",
						 "000001011001100111011010",
						 "000001011001100011011110",
						 "000001011001011111100010",
						 "000001011001011011100110",
						 "000001011001010111101010",
						 "000001011001010011101110",
						 "000001011001001111110010",
						 "000001011001001011110110",
						 "000001011001000111111010",
						 "000001011010000011001101",
						 "000001011001111111010000",
						 "000001011001111011010011",
						 "000001011001110111010110",
						 "000001011001110011011001",
						 "000001011001101111011100",
						 "000001011001101011011111",
						 "000001011001100111100010",
						 "000001011001100011100101",
						 "000001011001011111101000",
						 "000001011001011011101011",
						 "000001011001010111101110",
						 "000001011001010011110001",
						 "000001011001001111110100",
						 "000001011001001011110111",
						 "000001011001000111111010",
						 "000001011010000011001101",
						 "000001011001111111010000",
						 "000001011001111011010011",
						 "000001011001110111010110",
						 "000001011001110011011001",
						 "000001011001101111011100",
						 "000001011001101011011111",
						 "000001011001100111100010",
						 "000001011001100011100101",
						 "000001011001011111101000",
						 "000001011001011011101011",
						 "000001011001010111101110",
						 "000001011001010011110001",
						 "000001011001001111110100",
						 "000001011001001011110111",
						 "000001011001000111111010",
						 "000001010111100000001111",
						 "000001010111011100010010",
						 "000001010111011000010101",
						 "000001010111010100011000",
						 "000001010111010000011011",
						 "000001010111001100011110",
						 "000001010111001000100001",
						 "000001010111000100100100",
						 "000001010111000000100111",
						 "000001010110111100101010",
						 "000001010110111000101101",
						 "000001010110110100110000",
						 "000001010110110000110011",
						 "000001010110101100110110",
						 "000001010110101000111001",
						 "000001010110100100111100",
						 "000001010111100000001111",
						 "000001010111011100010010",
						 "000001010111011000010101",
						 "000001010111010100011000",
						 "000001010111010000011011",
						 "000001010111001100011110",
						 "000001010111001000100001",
						 "000001010111000100100100",
						 "000001010111000000100111",
						 "000001010110111100101010",
						 "000001010110111000101101",
						 "000001010110110100110000",
						 "000001010110110000110011",
						 "000001010110101100110110",
						 "000001010110101000111001",
						 "000001010110100100111100",
						 "000001010111100000001111",
						 "000001010111011100010010",
						 "000001010111011000010101",
						 "000001010111010100011000",
						 "000001010111010000011011",
						 "000001010111001100011110",
						 "000001010111001000100001",
						 "000001010111000100100100",
						 "000001010111000000100111",
						 "000001010110111100101010",
						 "000001010110111000101101",
						 "000001010110110100110000",
						 "000001010110110000110011",
						 "000001010110101100110110",
						 "000001010110101000111001",
						 "000001010110100100111100",
						 "000001010100111101010001",
						 "000001010100111001010100",
						 "000001010100110101010111",
						 "000001010100110001011010",
						 "000001010100101101011101",
						 "000001010100101001100000",
						 "000001010100100101100011",
						 "000001010100100001100110",
						 "000001010100011101101001",
						 "000001010100011001101100",
						 "000001010100010101101111",
						 "000001010100010001110010",
						 "000001010100001101110101",
						 "000001010100001001111000",
						 "000001010100000101111011",
						 "000001010100000001111110",
						 "000001010100111101010001",
						 "000001010100111001010100",
						 "000001010100110101010111",
						 "000001010100110001011010",
						 "000001010100101101011101",
						 "000001010100101001100000",
						 "000001010100100101100011",
						 "000001010100100001100110",
						 "000001010100011101101001",
						 "000001010100011001101100",
						 "000001010100010101101111",
						 "000001010100010001110010",
						 "000001010100001101110101",
						 "000001010100001001111000",
						 "000001010100000101111011",
						 "000001010100000001111110",
						 "000001010010011010010011",
						 "000001010010010110010110",
						 "000001010010010010011001",
						 "000001010010001110011100",
						 "000001010010001010011111",
						 "000001010010000110100010",
						 "000001010010000010100101",
						 "000001010001111110101000",
						 "000001010001111010101011",
						 "000001010001110110101110",
						 "000001010001110010110001",
						 "000001010001101110110100",
						 "000001010001101010110111",
						 "000001010001100110111010",
						 "000001010001100010111101",
						 "000001010001011111000000",
						 "000001010010011010010011",
						 "000001010010010110010110",
						 "000001010010010010011001",
						 "000001010010001110011100",
						 "000001010010001010011111",
						 "000001010010000110100010",
						 "000001010010000010100101",
						 "000001010001111110101000",
						 "000001010001111010101011",
						 "000001010001110110101110",
						 "000001010001110010110001",
						 "000001010001101110110100",
						 "000001010001101010110111",
						 "000001010001100110111010",
						 "000001010001100010111101",
						 "000001010001011111000000",
						 "000001010010011010010011",
						 "000001010010010110010110",
						 "000001010010010010011001",
						 "000001010010001110011100",
						 "000001010010001010011111",
						 "000001010010000110100010",
						 "000001010010000010100101",
						 "000001010001111110101000",
						 "000001010001111010101011",
						 "000001010001110110101110",
						 "000001010001110010110001",
						 "000001010001101110110100",
						 "000001010001101010110111",
						 "000001010001100110111010",
						 "000001010001100010111101",
						 "000001010001011111000000",
						 "000001001111110111010101",
						 "000001001111110011011000",
						 "000001001111101111011011",
						 "000001001111101011011110",
						 "000001001111100111100001",
						 "000001001111100011100100",
						 "000001001111011111100111",
						 "000001001111011011101010",
						 "000001001111010111101101",
						 "000001001111010011110000",
						 "000001001111001111110011",
						 "000001001111001011110110",
						 "000001001111000111111001",
						 "000001001111000011111100",
						 "000001001110111111111111",
						 "000001001110111100000010",
						 "000001001111110111010101",
						 "000001001111110011011000",
						 "000001001111101111011011",
						 "000001001111101011011110",
						 "000001001111100111100001",
						 "000001001111100011100100",
						 "000001001111011111100111",
						 "000001001111011011101010",
						 "000001001111010111101101",
						 "000001001111010011110000",
						 "000001001111001111110011",
						 "000001001111001011110110",
						 "000001001111000111111001",
						 "000001001111000011111100",
						 "000001001110111111111111",
						 "000001001110111100000010",
						 "000001001101010100010111",
						 "000001001101010000011010",
						 "000001001101001100011101",
						 "000001001101001000100000",
						 "000001001101000100100011",
						 "000001001101000000100110",
						 "000001001100111100101001",
						 "000001001100111000101100",
						 "000001001100110100101111",
						 "000001001100110000110010",
						 "000001001100101100110101",
						 "000001001100101000111000",
						 "000001001100100100111011",
						 "000001001100100000111110",
						 "000001001100011101000001",
						 "000001001100011001000100",
						 "000001001101010100010111",
						 "000001001101010000011010",
						 "000001001101001100011101",
						 "000001001101001000100000",
						 "000001001101000100100011",
						 "000001001101000000100110",
						 "000001001100111100101001",
						 "000001001100111000101100",
						 "000001001100110100101111",
						 "000001001100110000110010",
						 "000001001100101100110101",
						 "000001001100101000111000",
						 "000001001100100100111011",
						 "000001001100100000111110",
						 "000001001100011101000001",
						 "000001001100011001000100",
						 "000001001101010100010111",
						 "000001001101010000011010",
						 "000001001101001100011101",
						 "000001001101001000100000",
						 "000001001101000100100011",
						 "000001001101000000100110",
						 "000001001100111100101001",
						 "000001001100111000101100",
						 "000001001100110100101111",
						 "000001001100110000110010",
						 "000001001100101100110101",
						 "000001001100101000111000",
						 "000001001100100100111011",
						 "000001001100100000111110",
						 "000001001100011101000001",
						 "000001001100011001000100",
						 "000001001010110001011001",
						 "000001001010101101011100",
						 "000001001010101001011111",
						 "000001001010100101100010",
						 "000001001010100001100101",
						 "000001001010011101101000",
						 "000001001010011001101011",
						 "000001001010010101101110",
						 "000001001010010001110001",
						 "000001001010001101110100",
						 "000001001010001001110111",
						 "000001001010000101111010",
						 "000001001010000001111101",
						 "000001001001111110000000",
						 "000001001001111010000011",
						 "000001001001110110000110",
						 "000001001010110001011001",
						 "000001001010101101011100",
						 "000001001010101001011111",
						 "000001001010100101100010",
						 "000001001010100001100101",
						 "000001001010011101101000",
						 "000001001010011001101011",
						 "000001001010010101101110",
						 "000001001010010001110001",
						 "000001001010001101110100",
						 "000001001010001001110111",
						 "000001001010000101111010",
						 "000001001010000001111101",
						 "000001001001111110000000",
						 "000001001001111010000011",
						 "000001001001110110000110",
						 "000001001000001110011011",
						 "000001001000001010011110",
						 "000001001000000110100001",
						 "000001001000000010100100",
						 "000001000111111110100111",
						 "000001000111111010101010",
						 "000001000111110110101101",
						 "000001000111110010110000",
						 "000001000111101110110011",
						 "000001000111101010110110",
						 "000001000111100110111001",
						 "000001000111100010111100",
						 "000001000111011110111111",
						 "000001000111011011000010",
						 "000001000111010111000101",
						 "000001000111010011001000",
						 "000001001000001110011011",
						 "000001001000001010011110",
						 "000001001000000110100001",
						 "000001001000000010100100",
						 "000001000111111110100111",
						 "000001000111111010101010",
						 "000001000111110110101101",
						 "000001000111110010110000",
						 "000001000111101110110011",
						 "000001000111101010110110",
						 "000001000111100110111001",
						 "000001000111100010111100",
						 "000001000111011110111111",
						 "000001000111011011000010",
						 "000001000111010111000101",
						 "000001000111010011001000",
						 "000001001000001110011011",
						 "000001001000001010011110",
						 "000001001000000110100001",
						 "000001001000000010100100",
						 "000001000111111110100111",
						 "000001000111111010101010",
						 "000001000111110110101101",
						 "000001000111110010110000",
						 "000001000111101110110011",
						 "000001000111101010110110",
						 "000001000111100110111001",
						 "000001000111100010111100",
						 "000001000111011110111111",
						 "000001000111011011000010",
						 "000001000111010111000101",
						 "000001000111010011001000",
						 "000001000101101011101100",
						 "000001000101100111101110",
						 "000001000101100011110000",
						 "000001000101011111110010",
						 "000001000101011011110100",
						 "000001000101010111110110",
						 "000001000101010011111000",
						 "000001000101001111111010",
						 "000001000101001011111100",
						 "000001000101000111111110",
						 "000001000101000100000000",
						 "000001000101000000000010",
						 "000001000100111100000100",
						 "000001000100111000000110",
						 "000001000100110100001000",
						 "000001000100110000001010",
						 "000001000101101011101100",
						 "000001000101100111101110",
						 "000001000101100011110000",
						 "000001000101011111110010",
						 "000001000101011011110100",
						 "000001000101010111110110",
						 "000001000101010011111000",
						 "000001000101001111111010",
						 "000001000101001011111100",
						 "000001000101000111111110",
						 "000001000101000100000000",
						 "000001000101000000000010",
						 "000001000100111100000100",
						 "000001000100111000000110",
						 "000001000100110100001000",
						 "000001000100110000001010",
						 "000001000101101011101100",
						 "000001000101100111101110",
						 "000001000101100011110000",
						 "000001000101011111110010",
						 "000001000101011011110100",
						 "000001000101010111110110",
						 "000001000101010011111000",
						 "000001000101001111111010",
						 "000001000101001011111100",
						 "000001000101000111111110",
						 "000001000101000100000000",
						 "000001000101000000000010",
						 "000001000100111100000100",
						 "000001000100111000000110",
						 "000001000100110100001000",
						 "000001000100110000001010",
						 "000001000011001000101110",
						 "000001000011000100110000",
						 "000001000011000000110010",
						 "000001000010111100110100",
						 "000001000010111000110110",
						 "000001000010110100111000",
						 "000001000010110000111010",
						 "000001000010101100111100",
						 "000001000010101000111110",
						 "000001000010100101000000",
						 "000001000010100001000010",
						 "000001000010011101000100",
						 "000001000010011001000110",
						 "000001000010010101001000",
						 "000001000010010001001010",
						 "000001000010001101001100",
						 "000001000011001000101110",
						 "000001000011000100110000",
						 "000001000011000000110010",
						 "000001000010111100110100",
						 "000001000010111000110110",
						 "000001000010110100111000",
						 "000001000010110000111010",
						 "000001000010101100111100",
						 "000001000010101000111110",
						 "000001000010100101000000",
						 "000001000010100001000010",
						 "000001000010011101000100",
						 "000001000010011001000110",
						 "000001000010010101001000",
						 "000001000010010001001010",
						 "000001000010001101001100",
						 "000001000000100101110000",
						 "000001000000100001110010",
						 "000001000000011101110100",
						 "000001000000011001110110",
						 "000001000000010101111000",
						 "000001000000010001111010",
						 "000001000000001101111100",
						 "000001000000001001111110",
						 "000001000000000110000000",
						 "000001000000000010000010",
						 "000000111111111110000100",
						 "000000111111111010000110",
						 "000000111111110110001000",
						 "000000111111110010001010",
						 "000000111111101110001100",
						 "000000111111101010001110",
						 "000001000000100101110000",
						 "000001000000100001110010",
						 "000001000000011101110100",
						 "000001000000011001110110",
						 "000001000000010101111000",
						 "000001000000010001111010",
						 "000001000000001101111100",
						 "000001000000001001111110",
						 "000001000000000110000000",
						 "000001000000000010000010",
						 "000000111111111110000100",
						 "000000111111111010000110",
						 "000000111111110110001000",
						 "000000111111110010001010",
						 "000000111111101110001100",
						 "000000111111101010001110",
						 "000001000000100101110000",
						 "000001000000100001110010",
						 "000001000000011101110100",
						 "000001000000011001110110",
						 "000001000000010101111000",
						 "000001000000010001111010",
						 "000001000000001101111100",
						 "000001000000001001111110",
						 "000001000000000110000000",
						 "000001000000000010000010",
						 "000000111111111110000100",
						 "000000111111111010000110",
						 "000000111111110110001000",
						 "000000111111110010001010",
						 "000000111111101110001100",
						 "000000111111101010001110",
						 "000000111110000010110010",
						 "000000111101111110110100",
						 "000000111101111010110110",
						 "000000111101110110111000",
						 "000000111101110010111010",
						 "000000111101101110111100",
						 "000000111101101010111110",
						 "000000111101100111000000",
						 "000000111101100011000010",
						 "000000111101011111000100",
						 "000000111101011011000110",
						 "000000111101010111001000",
						 "000000111101010011001010",
						 "000000111101001111001100",
						 "000000111101001011001110",
						 "000000111101000111010000",
						 "000000111110000010110010",
						 "000000111101111110110100",
						 "000000111101111010110110",
						 "000000111101110110111000",
						 "000000111101110010111010",
						 "000000111101101110111100",
						 "000000111101101010111110",
						 "000000111101100111000000",
						 "000000111101100011000010",
						 "000000111101011111000100",
						 "000000111101011011000110",
						 "000000111101010111001000",
						 "000000111101010011001010",
						 "000000111101001111001100",
						 "000000111101001011001110",
						 "000000111101000111010000",
						 "000000111011011111110100",
						 "000000111011011011110110",
						 "000000111011010111111000",
						 "000000111011010011111010",
						 "000000111011001111111100",
						 "000000111011001011111110",
						 "000000111011001000000000",
						 "000000111011000100000010",
						 "000000111011000000000100",
						 "000000111010111100000110",
						 "000000111010111000001000",
						 "000000111010110100001010",
						 "000000111010110000001100",
						 "000000111010101100001110",
						 "000000111010101000010000",
						 "000000111010100100010010",
						 "000000111011011111110100",
						 "000000111011011011110110",
						 "000000111011010111111000",
						 "000000111011010011111010",
						 "000000111011001111111100",
						 "000000111011001011111110",
						 "000000111011001000000000",
						 "000000111011000100000010",
						 "000000111011000000000100",
						 "000000111010111100000110",
						 "000000111010111000001000",
						 "000000111010110100001010",
						 "000000111010110000001100",
						 "000000111010101100001110",
						 "000000111010101000010000",
						 "000000111010100100010010",
						 "000000111011011111110100",
						 "000000111011011011110110",
						 "000000111011010111111000",
						 "000000111011010011111010",
						 "000000111011001111111100",
						 "000000111011001011111110",
						 "000000111011001000000000",
						 "000000111011000100000010",
						 "000000111011000000000100",
						 "000000111010111100000110",
						 "000000111010111000001000",
						 "000000111010110100001010",
						 "000000111010110000001100",
						 "000000111010101100001110",
						 "000000111010101000010000",
						 "000000111010100100010010",
						 "000000111000111100110110",
						 "000000111000111000111000",
						 "000000111000110100111010",
						 "000000111000110000111100",
						 "000000111000101100111110",
						 "000000111000101001000000",
						 "000000111000100101000010",
						 "000000111000100001000100",
						 "000000111000011101000110",
						 "000000111000011001001000",
						 "000000111000010101001010",
						 "000000111000010001001100",
						 "000000111000001101001110",
						 "000000111000001001010000",
						 "000000111000000101010010",
						 "000000111000000001010100",
						 "000000111000111100110110",
						 "000000111000111000111000",
						 "000000111000110100111010",
						 "000000111000110000111100",
						 "000000111000101100111110",
						 "000000111000101001000000",
						 "000000111000100101000010",
						 "000000111000100001000100",
						 "000000111000011101000110",
						 "000000111000011001001000",
						 "000000111000010101001010",
						 "000000111000010001001100",
						 "000000111000001101001110",
						 "000000111000001001010000",
						 "000000111000000101010010",
						 "000000111000000001010100",
						 "000000110110011001111000",
						 "000000110110010101111010",
						 "000000110110010001111100",
						 "000000110110001101111110",
						 "000000110110001010000000",
						 "000000110110000110000010",
						 "000000110110000010000100",
						 "000000110101111110000110",
						 "000000110101111010001000",
						 "000000110101110110001010",
						 "000000110101110010001100",
						 "000000110101101110001110",
						 "000000110101101010010000",
						 "000000110101100110010010",
						 "000000110101100010010100",
						 "000000110101011110010110",
						 "000000110110011001111000",
						 "000000110110010101111010",
						 "000000110110010001111100",
						 "000000110110001101111110",
						 "000000110110001010000000",
						 "000000110110000110000010",
						 "000000110110000010000100",
						 "000000110101111110000110",
						 "000000110101111010001000",
						 "000000110101110110001010",
						 "000000110101110010001100",
						 "000000110101101110001110",
						 "000000110101101010010000",
						 "000000110101100110010010",
						 "000000110101100010010100",
						 "000000110101011110010110",
						 "000000110110011001111000",
						 "000000110110010101111010",
						 "000000110110010001111100",
						 "000000110110001101111110",
						 "000000110110001010000000",
						 "000000110110000110000010",
						 "000000110110000010000100",
						 "000000110101111110000110",
						 "000000110101111010001000",
						 "000000110101110110001010",
						 "000000110101110010001100",
						 "000000110101101110001110",
						 "000000110101101010010000",
						 "000000110101100110010010",
						 "000000110101100010010100",
						 "000000110101011110010110",
						 "000000110011110110111010",
						 "000000110011110010111100",
						 "000000110011101110111110",
						 "000000110011101011000000",
						 "000000110011100111000010",
						 "000000110011100011000100",
						 "000000110011011111000110",
						 "000000110011011011001000",
						 "000000110011010111001010",
						 "000000110011010011001100",
						 "000000110011001111001110",
						 "000000110011001011010000",
						 "000000110011000111010010",
						 "000000110011000011010100",
						 "000000110010111111010110",
						 "000000110010111011011000",
						 "000000110011110110111010",
						 "000000110011110010111100",
						 "000000110011101110111110",
						 "000000110011101011000000",
						 "000000110011100111000010",
						 "000000110011100011000100",
						 "000000110011011111000110",
						 "000000110011011011001000",
						 "000000110011010111001010",
						 "000000110011010011001100",
						 "000000110011001111001110",
						 "000000110011001011010000",
						 "000000110011000111010010",
						 "000000110011000011010100",
						 "000000110010111111010110",
						 "000000110010111011011000",
						 "000000110011110110111010",
						 "000000110011110010111100",
						 "000000110011101110111110",
						 "000000110011101011000000",
						 "000000110011100111000010",
						 "000000110011100011000100",
						 "000000110011011111000110",
						 "000000110011011011001000",
						 "000000110011010111001010",
						 "000000110011010011001100",
						 "000000110011001111001110",
						 "000000110011001011010000",
						 "000000110011000111010010",
						 "000000110011000011010100",
						 "000000110010111111010110",
						 "000000110010111011011000",
						 "000000110001010011111100",
						 "000000110001001111111110",
						 "000000110001001100000000",
						 "000000110001001000000010",
						 "000000110001000100000100",
						 "000000110001000000000110",
						 "000000110000111100001000",
						 "000000110000111000001010",
						 "000000110000110100001100",
						 "000000110000110000001110",
						 "000000110000101100010000",
						 "000000110000101000010010",
						 "000000110000100100010100",
						 "000000110000100000010110",
						 "000000110000011100011000",
						 "000000110000011000011010",
						 "000000110001010011111100",
						 "000000110001001111111110",
						 "000000110001001100000000",
						 "000000110001001000000010",
						 "000000110001000100000100",
						 "000000110001000000000110",
						 "000000110000111100001000",
						 "000000110000111000001010",
						 "000000110000110100001100",
						 "000000110000110000001110",
						 "000000110000101100010000",
						 "000000110000101000010010",
						 "000000110000100100010100",
						 "000000110000100000010110",
						 "000000110000011100011000",
						 "000000110000011000011010",
						 "000000101110110000111110",
						 "000000101110101101000000",
						 "000000101110101001000010",
						 "000000101110100101000100",
						 "000000101110100001000110",
						 "000000101110011101001000",
						 "000000101110011001001010",
						 "000000101110010101001100",
						 "000000101110010001001110",
						 "000000101110001101010000",
						 "000000101110001001010010",
						 "000000101110000101010100",
						 "000000101110000001010110",
						 "000000101101111101011000",
						 "000000101101111001011010",
						 "000000101101110101011100",
						 "000000101110110000111110",
						 "000000101110101101000000",
						 "000000101110101001000010",
						 "000000101110100101000100",
						 "000000101110100001000110",
						 "000000101110011101001000",
						 "000000101110011001001010",
						 "000000101110010101001100",
						 "000000101110010001001110",
						 "000000101110001101010000",
						 "000000101110001001010010",
						 "000000101110000101010100",
						 "000000101110000001010110",
						 "000000101101111101011000",
						 "000000101101111001011010",
						 "000000101101110101011100",
						 "000000101110110000111110",
						 "000000101110101101000000",
						 "000000101110101001000010",
						 "000000101110100101000100",
						 "000000101110100001000110",
						 "000000101110011101001000",
						 "000000101110011001001010",
						 "000000101110010101001100",
						 "000000101110010001001110",
						 "000000101110001101010000",
						 "000000101110001001010010",
						 "000000101110000101010100",
						 "000000101110000001010110",
						 "000000101101111101011000",
						 "000000101101111001011010",
						 "000000101101110101011100",
						 "000000101100001110000000",
						 "000000101100001010000010",
						 "000000101100000110000100",
						 "000000101100000010000110",
						 "000000101011111110001000",
						 "000000101011111010001010",
						 "000000101011110110001100",
						 "000000101011110010001110",
						 "000000101011101110010000",
						 "000000101011101010010010",
						 "000000101011100110010100",
						 "000000101011100010010110",
						 "000000101011011110011000",
						 "000000101011011010011010",
						 "000000101011010110011100",
						 "000000101011010010011110",
						 "000000101100001110000000",
						 "000000101100001010000010",
						 "000000101100000110000100",
						 "000000101100000010000110",
						 "000000101011111110001000",
						 "000000101011111010001010",
						 "000000101011110110001100",
						 "000000101011110010001110",
						 "000000101011101110010000",
						 "000000101011101010010010",
						 "000000101011100110010100",
						 "000000101011100010010110",
						 "000000101011011110011000",
						 "000000101011011010011010",
						 "000000101011010110011100",
						 "000000101011010010011110",
						 "000000101001101011000010",
						 "000000101001100111000100",
						 "000000101001100011000110",
						 "000000101001011111001000",
						 "000000101001011011001010",
						 "000000101001010111001100",
						 "000000101001010011001110",
						 "000000101001001111010000",
						 "000000101001001011010010",
						 "000000101001000111010100",
						 "000000101001000011010110",
						 "000000101000111111011000",
						 "000000101000111011011010",
						 "000000101000110111011100",
						 "000000101000110011011110",
						 "000000101000101111100000",
						 "000000101001101011000010",
						 "000000101001100111000100",
						 "000000101001100011000110",
						 "000000101001011111001000",
						 "000000101001011011001010",
						 "000000101001010111001100",
						 "000000101001010011001110",
						 "000000101001001111010000",
						 "000000101001001011010010",
						 "000000101001000111010100",
						 "000000101001000011010110",
						 "000000101000111111011000",
						 "000000101000111011011010",
						 "000000101000110111011100",
						 "000000101000110011011110",
						 "000000101000101111100000",
						 "000000101001101011010001",
						 "000000101001100111010010",
						 "000000101001100011010011",
						 "000000101001011111010100",
						 "000000101001011011010101",
						 "000000101001010111010110",
						 "000000101001010011010111",
						 "000000101001001111011000",
						 "000000101001001011011001",
						 "000000101001000111011010",
						 "000000101001000011011011",
						 "000000101000111111011100",
						 "000000101000111011011101",
						 "000000101000110111011110",
						 "000000101000110011011111",
						 "000000101000101111100000",
						 "000000100111001000010011",
						 "000000100111000100010100",
						 "000000100111000000010101",
						 "000000100110111100010110",
						 "000000100110111000010111",
						 "000000100110110100011000",
						 "000000100110110000011001",
						 "000000100110101100011010",
						 "000000100110101000011011",
						 "000000100110100100011100",
						 "000000100110100000011101",
						 "000000100110011100011110",
						 "000000100110011000011111",
						 "000000100110010100100000",
						 "000000100110010000100001",
						 "000000100110001100100010",
						 "000000100111001000010011",
						 "000000100111000100010100",
						 "000000100111000000010101",
						 "000000100110111100010110",
						 "000000100110111000010111",
						 "000000100110110100011000",
						 "000000100110110000011001",
						 "000000100110101100011010",
						 "000000100110101000011011",
						 "000000100110100100011100",
						 "000000100110100000011101",
						 "000000100110011100011110",
						 "000000100110011000011111",
						 "000000100110010100100000",
						 "000000100110010000100001",
						 "000000100110001100100010",
						 "000000100100100101010101",
						 "000000100100100001010110",
						 "000000100100011101010111",
						 "000000100100011001011000",
						 "000000100100010101011001",
						 "000000100100010001011010",
						 "000000100100001101011011",
						 "000000100100001001011100",
						 "000000100100000101011101",
						 "000000100100000001011110",
						 "000000100011111101011111",
						 "000000100011111001100000",
						 "000000100011110101100001",
						 "000000100011110001100010",
						 "000000100011101101100011",
						 "000000100011101001100100",
						 "000000100100100101010101",
						 "000000100100100001010110",
						 "000000100100011101010111",
						 "000000100100011001011000",
						 "000000100100010101011001",
						 "000000100100010001011010",
						 "000000100100001101011011",
						 "000000100100001001011100",
						 "000000100100000101011101",
						 "000000100100000001011110",
						 "000000100011111101011111",
						 "000000100011111001100000",
						 "000000100011110101100001",
						 "000000100011110001100010",
						 "000000100011101101100011",
						 "000000100011101001100100",
						 "000000100100100101010101",
						 "000000100100100001010110",
						 "000000100100011101010111",
						 "000000100100011001011000",
						 "000000100100010101011001",
						 "000000100100010001011010",
						 "000000100100001101011011",
						 "000000100100001001011100",
						 "000000100100000101011101",
						 "000000100100000001011110",
						 "000000100011111101011111",
						 "000000100011111001100000",
						 "000000100011110101100001",
						 "000000100011110001100010",
						 "000000100011101101100011",
						 "000000100011101001100100",
						 "000000100010000010010111",
						 "000000100001111110011000",
						 "000000100001111010011001",
						 "000000100001110110011010",
						 "000000100001110010011011",
						 "000000100001101110011100",
						 "000000100001101010011101",
						 "000000100001100110011110",
						 "000000100001100010011111",
						 "000000100001011110100000",
						 "000000100001011010100001",
						 "000000100001010110100010",
						 "000000100001010010100011",
						 "000000100001001110100100",
						 "000000100001001010100101",
						 "000000100001000110100110",
						 "000000100010000010010111",
						 "000000100001111110011000",
						 "000000100001111010011001",
						 "000000100001110110011010",
						 "000000100001110010011011",
						 "000000100001101110011100",
						 "000000100001101010011101",
						 "000000100001100110011110",
						 "000000100001100010011111",
						 "000000100001011110100000",
						 "000000100001011010100001",
						 "000000100001010110100010",
						 "000000100001010010100011",
						 "000000100001001110100100",
						 "000000100001001010100101",
						 "000000100001000110100110",
						 "000000100010000010010111",
						 "000000100001111110011000",
						 "000000100001111010011001",
						 "000000100001110110011010",
						 "000000100001110010011011",
						 "000000100001101110011100",
						 "000000100001101010011101",
						 "000000100001100110011110",
						 "000000100001100010011111",
						 "000000100001011110100000",
						 "000000100001011010100001",
						 "000000100001010110100010",
						 "000000100001010010100011",
						 "000000100001001110100100",
						 "000000100001001010100101",
						 "000000100001000110100110",
						 "000000011111011111011001",
						 "000000011111011011011010",
						 "000000011111010111011011",
						 "000000011111010011011100",
						 "000000011111001111011101",
						 "000000011111001011011110",
						 "000000011111000111011111",
						 "000000011111000011100000",
						 "000000011110111111100001",
						 "000000011110111011100010",
						 "000000011110110111100011",
						 "000000011110110011100100",
						 "000000011110101111100101",
						 "000000011110101011100110",
						 "000000011110100111100111",
						 "000000011110100011101000",
						 "000000011111011111011001",
						 "000000011111011011011010",
						 "000000011111010111011011",
						 "000000011111010011011100",
						 "000000011111001111011101",
						 "000000011111001011011110",
						 "000000011111000111011111",
						 "000000011111000011100000",
						 "000000011110111111100001",
						 "000000011110111011100010",
						 "000000011110110111100011",
						 "000000011110110011100100",
						 "000000011110101111100101",
						 "000000011110101011100110",
						 "000000011110100111100111",
						 "000000011110100011101000",
						 "000000011100111100011011",
						 "000000011100111000011100",
						 "000000011100110100011101",
						 "000000011100110000011110",
						 "000000011100101100011111",
						 "000000011100101000100000",
						 "000000011100100100100001",
						 "000000011100100000100010",
						 "000000011100011100100011",
						 "000000011100011000100100",
						 "000000011100010100100101",
						 "000000011100010000100110",
						 "000000011100001100100111",
						 "000000011100001000101000",
						 "000000011100000100101001",
						 "000000011100000000101010",
						 "000000011100111100011011",
						 "000000011100111000011100",
						 "000000011100110100011101",
						 "000000011100110000011110",
						 "000000011100101100011111",
						 "000000011100101000100000",
						 "000000011100100100100001",
						 "000000011100100000100010",
						 "000000011100011100100011",
						 "000000011100011000100100",
						 "000000011100010100100101",
						 "000000011100010000100110",
						 "000000011100001100100111",
						 "000000011100001000101000",
						 "000000011100000100101001",
						 "000000011100000000101010",
						 "000000011100111100011011",
						 "000000011100111000011100",
						 "000000011100110100011101",
						 "000000011100110000011110",
						 "000000011100101100011111",
						 "000000011100101000100000",
						 "000000011100100100100001",
						 "000000011100100000100010",
						 "000000011100011100100011",
						 "000000011100011000100100",
						 "000000011100010100100101",
						 "000000011100010000100110",
						 "000000011100001100100111",
						 "000000011100001000101000",
						 "000000011100000100101001",
						 "000000011100000000101010",
						 "000000011010011001011101",
						 "000000011010010101011110",
						 "000000011010010001011111",
						 "000000011010001101100000",
						 "000000011010001001100001",
						 "000000011010000101100010",
						 "000000011010000001100011",
						 "000000011001111101100100",
						 "000000011001111001100101",
						 "000000011001110101100110",
						 "000000011001110001100111",
						 "000000011001101101101000",
						 "000000011001101001101001",
						 "000000011001100101101010",
						 "000000011001100001101011",
						 "000000011001011101101100",
						 "000000011010011001011101",
						 "000000011010010101011110",
						 "000000011010010001011111",
						 "000000011010001101100000",
						 "000000011010001001100001",
						 "000000011010000101100010",
						 "000000011010000001100011",
						 "000000011001111101100100",
						 "000000011001111001100101",
						 "000000011001110101100110",
						 "000000011001110001100111",
						 "000000011001101101101000",
						 "000000011001101001101001",
						 "000000011001100101101010",
						 "000000011001100001101011",
						 "000000011001011101101100",
						 "000000010111110110011111",
						 "000000010111110010100000",
						 "000000010111101110100001",
						 "000000010111101010100010",
						 "000000010111100110100011",
						 "000000010111100010100100",
						 "000000010111011110100101",
						 "000000010111011010100110",
						 "000000010111010110100111",
						 "000000010111010010101000",
						 "000000010111001110101001",
						 "000000010111001010101010",
						 "000000010111000110101011",
						 "000000010111000010101100",
						 "000000010110111110101101",
						 "000000010110111010101110",
						 "000000010111110110011111",
						 "000000010111110010100000",
						 "000000010111101110100001",
						 "000000010111101010100010",
						 "000000010111100110100011",
						 "000000010111100010100100",
						 "000000010111011110100101",
						 "000000010111011010100110",
						 "000000010111010110100111",
						 "000000010111010010101000",
						 "000000010111001110101001",
						 "000000010111001010101010",
						 "000000010111000110101011",
						 "000000010111000010101100",
						 "000000010110111110101101",
						 "000000010110111010101110",
						 "000000010111110110011111",
						 "000000010111110010100000",
						 "000000010111101110100001",
						 "000000010111101010100010",
						 "000000010111100110100011",
						 "000000010111100010100100",
						 "000000010111011110100101",
						 "000000010111011010100110",
						 "000000010111010110100111",
						 "000000010111010010101000",
						 "000000010111001110101001",
						 "000000010111001010101010",
						 "000000010111000110101011",
						 "000000010111000010101100",
						 "000000010110111110101101",
						 "000000010110111010101110",
						 "000000010101010011100001",
						 "000000010101001111100010",
						 "000000010101001011100011",
						 "000000010101000111100100",
						 "000000010101000011100101",
						 "000000010100111111100110",
						 "000000010100111011100111",
						 "000000010100110111101000",
						 "000000010100110011101001",
						 "000000010100101111101010",
						 "000000010100101011101011",
						 "000000010100100111101100",
						 "000000010100100011101101",
						 "000000010100011111101110",
						 "000000010100011011101111",
						 "000000010100010111110000",
						 "000000010101010011100001",
						 "000000010101001111100010",
						 "000000010101001011100011",
						 "000000010101000111100100",
						 "000000010101000011100101",
						 "000000010100111111100110",
						 "000000010100111011100111",
						 "000000010100110111101000",
						 "000000010100110011101001",
						 "000000010100101111101010",
						 "000000010100101011101011",
						 "000000010100100111101100",
						 "000000010100100011101101",
						 "000000010100011111101110",
						 "000000010100011011101111",
						 "000000010100010111110000",
						 "000000010010110000100011",
						 "000000010010101100100100",
						 "000000010010101000100101",
						 "000000010010100100100110",
						 "000000010010100000100111",
						 "000000010010011100101000",
						 "000000010010011000101001",
						 "000000010010010100101010",
						 "000000010010010000101011",
						 "000000010010001100101100",
						 "000000010010001000101101",
						 "000000010010000100101110",
						 "000000010010000000101111",
						 "000000010001111100110000",
						 "000000010001111000110001",
						 "000000010001110100110010",
						 "000000010010110000100011",
						 "000000010010101100100100",
						 "000000010010101000100101",
						 "000000010010100100100110",
						 "000000010010100000100111",
						 "000000010010011100101000",
						 "000000010010011000101001",
						 "000000010010010100101010",
						 "000000010010010000101011",
						 "000000010010001100101100",
						 "000000010010001000101101",
						 "000000010010000100101110",
						 "000000010010000000101111",
						 "000000010001111100110000",
						 "000000010001111000110001",
						 "000000010001110100110010",
						 "000000010010110000100011",
						 "000000010010101100100100",
						 "000000010010101000100101",
						 "000000010010100100100110",
						 "000000010010100000100111",
						 "000000010010011100101000",
						 "000000010010011000101001",
						 "000000010010010100101010",
						 "000000010010010000101011",
						 "000000010010001100101100",
						 "000000010010001000101101",
						 "000000010010000100101110",
						 "000000010010000000101111",
						 "000000010001111100110000",
						 "000000010001111000110001",
						 "000000010001110100110010",
						 "000000010000001101100101",
						 "000000010000001001100110",
						 "000000010000000101100111",
						 "000000010000000001101000",
						 "000000001111111101101001",
						 "000000001111111001101010",
						 "000000001111110101101011",
						 "000000001111110001101100",
						 "000000001111101101101101",
						 "000000001111101001101110",
						 "000000001111100101101111",
						 "000000001111100001110000",
						 "000000001111011101110001",
						 "000000001111011001110010",
						 "000000001111010101110011",
						 "000000001111010001110100",
						 "000000010000001101100101",
						 "000000010000001001100110",
						 "000000010000000101100111",
						 "000000010000000001101000",
						 "000000001111111101101001",
						 "000000001111111001101010",
						 "000000001111110101101011",
						 "000000001111110001101100",
						 "000000001111101101101101",
						 "000000001111101001101110",
						 "000000001111100101101111",
						 "000000001111100001110000",
						 "000000001111011101110001",
						 "000000001111011001110010",
						 "000000001111010101110011",
						 "000000001111010001110100",
						 "000000001101101010100111",
						 "000000001101100110101000",
						 "000000001101100010101001",
						 "000000001101011110101010",
						 "000000001101011010101011",
						 "000000001101010110101100",
						 "000000001101010010101101",
						 "000000001101001110101110",
						 "000000001101001010101111",
						 "000000001101000110110000",
						 "000000001101000010110001",
						 "000000001100111110110010",
						 "000000001100111010110011",
						 "000000001100110110110100",
						 "000000001100110010110101",
						 "000000001100101110110110",
						 "000000001101101010100111",
						 "000000001101100110101000",
						 "000000001101100010101001",
						 "000000001101011110101010",
						 "000000001101011010101011",
						 "000000001101010110101100",
						 "000000001101010010101101",
						 "000000001101001110101110",
						 "000000001101001010101111",
						 "000000001101000110110000",
						 "000000001101000010110001",
						 "000000001100111110110010",
						 "000000001100111010110011",
						 "000000001100110110110100",
						 "000000001100110010110101",
						 "000000001100101110110110",
						 "000000001101101010100111",
						 "000000001101100110101000",
						 "000000001101100010101001",
						 "000000001101011110101010",
						 "000000001101011010101011",
						 "000000001101010110101100",
						 "000000001101010010101101",
						 "000000001101001110101110",
						 "000000001101001010101111",
						 "000000001101000110110000",
						 "000000001101000010110001",
						 "000000001100111110110010",
						 "000000001100111010110011",
						 "000000001100110110110100",
						 "000000001100110010110101",
						 "000000001100101110110110",
						 "000000001011000111101001",
						 "000000001011000011101010",
						 "000000001010111111101011",
						 "000000001010111011101100",
						 "000000001010110111101101",
						 "000000001010110011101110",
						 "000000001010101111101111",
						 "000000001010101011110000",
						 "000000001010100111110001",
						 "000000001010100011110010",
						 "000000001010011111110011",
						 "000000001010011011110100",
						 "000000001010010111110101",
						 "000000001010010011110110",
						 "000000001010001111110111",
						 "000000001010001011111000",
						 "000000001011000111101001",
						 "000000001011000011101010",
						 "000000001010111111101011",
						 "000000001010111011101100",
						 "000000001010110111101101",
						 "000000001010110011101110",
						 "000000001010101111101111",
						 "000000001010101011110000",
						 "000000001010100111110001",
						 "000000001010100011110010",
						 "000000001010011111110011",
						 "000000001010011011110100",
						 "000000001010010111110101",
						 "000000001010010011110110",
						 "000000001010001111110111",
						 "000000001010001011111000",
						 "000000001011000111101001",
						 "000000001011000011101010",
						 "000000001010111111101011",
						 "000000001010111011101100",
						 "000000001010110111101101",
						 "000000001010110011101110",
						 "000000001010101111101111",
						 "000000001010101011110000",
						 "000000001010100111110001",
						 "000000001010100011110010",
						 "000000001010011111110011",
						 "000000001010011011110100",
						 "000000001010010111110101",
						 "000000001010010011110110",
						 "000000001010001111110111",
						 "000000001010001011111000",
						 "000000001000100100101011",
						 "000000001000100000101100",
						 "000000001000011100101101",
						 "000000001000011000101110",
						 "000000001000010100101111",
						 "000000001000010000110000",
						 "000000001000001100110001",
						 "000000001000001000110010",
						 "000000001000000100110011",
						 "000000001000000000110100",
						 "000000000111111100110101",
						 "000000000111111000110110",
						 "000000000111110100110111",
						 "000000000111110000111000",
						 "000000000111101100111001",
						 "000000000111101000111010",
						 "000000001000100100101011",
						 "000000001000100000101100",
						 "000000001000011100101101",
						 "000000001000011000101110",
						 "000000001000010100101111",
						 "000000001000010000110000",
						 "000000001000001100110001",
						 "000000001000001000110010",
						 "000000001000000100110011",
						 "000000001000000000110100",
						 "000000000111111100110101",
						 "000000000111111000110110",
						 "000000000111110100110111",
						 "000000000111110000111000",
						 "000000000111101100111001",
						 "000000000111101000111010",
						 "000000000110000001101101",
						 "000000000101111101101110",
						 "000000000101111001101111",
						 "000000000101110101110000",
						 "000000000101110001110001",
						 "000000000101101101110010",
						 "000000000101101001110011",
						 "000000000101100101110100",
						 "000000000101100001110101",
						 "000000000101011101110110",
						 "000000000101011001110111",
						 "000000000101010101111000",
						 "000000000101010001111001",
						 "000000000101001101111010",
						 "000000000101001001111011",
						 "000000000101000101111100",
						 "000000000110000001101101",
						 "000000000101111101101110",
						 "000000000101111001101111",
						 "000000000101110101110000",
						 "000000000101110001110001",
						 "000000000101101101110010",
						 "000000000101101001110011",
						 "000000000101100101110100",
						 "000000000101100001110101",
						 "000000000101011101110110",
						 "000000000101011001110111",
						 "000000000101010101111000",
						 "000000000101010001111001",
						 "000000000101001101111010",
						 "000000000101001001111011",
						 "000000000101000101111100",
						 "000000000110000001101101",
						 "000000000101111101101110",
						 "000000000101111001101111",
						 "000000000101110101110000",
						 "000000000101110001110001",
						 "000000000101101101110010",
						 "000000000101101001110011",
						 "000000000101100101110100",
						 "000000000101100001110101",
						 "000000000101011101110110",
						 "000000000101011001110111",
						 "000000000101010101111000",
						 "000000000101010001111001",
						 "000000000101001101111010",
						 "000000000101001001111011",
						 "000000000101000101111100",
						 "000000000011011110101111",
						 "000000000011011010110000",
						 "000000000011010110110001",
						 "000000000011010010110010",
						 "000000000011001110110011",
						 "000000000011001010110100",
						 "000000000011000110110101",
						 "000000000011000010110110",
						 "000000000010111110110111",
						 "000000000010111010111000",
						 "000000000010110110111001",
						 "000000000010110010111010",
						 "000000000010101110111011",
						 "000000000010101010111100",
						 "000000000010100110111101",
						 "000000000010100010111110",
						 "000000000011011110101111",
						 "000000000011011010110000",
						 "000000000011010110110001",
						 "000000000011010010110010",
						 "000000000011001110110011",
						 "000000000011001010110100",
						 "000000000011000110110101",
						 "000000000011000010110110",
						 "000000000010111110110111",
						 "000000000010111010111000",
						 "000000000010110110111001",
						 "000000000010110010111010",
						 "000000000010101110111011",
						 "000000000010101010111100",
						 "000000000010100110111101",
						 "000000000010100010111110",
						 "000000000000111011110001",
						 "000000000000110111110010",
						 "000000000000110011110011",
						 "000000000000101111110100",
						 "000000000000101011110101",
						 "000000000000100111110110",
						 "000000000000100011110111",
						 "000000000000011111111000",
						 "000000000000011011111001",
						 "000000000000010111111010",
						 "000000000000010011111011",
						 "000000000000001111111100",
						 "000000000000001011111101",
						 "000000000000000111111110",
						 "000000000000000011111111",
						 "000000000000000000000000",
						 "000000000000111011110001",
						 "000000000000110111110010",
						 "000000000000110011110011",
						 "000000000000101111110100",
						 "000000000000101011110101",
						 "000000000000100111110110",
						 "000000000000100011110111",
						 "000000000000011111111000",
						 "000000000000011011111001",
						 "000000000000010111111010",
						 "000000000000010011111011",
						 "000000000000001111111100",
						 "000000000000001011111101",
						 "000000000000000111111110",
						 "000000000000000011111111",
						 "000000000000000000000000",
						 "100000000000000000000000",
						 "100000000000000011111111",
						 "100000000000000111111110",
						 "100000000000001011111101",
						 "100000000000001111111100",
						 "100000000000010011111011",
						 "100000000000010111111010",
						 "100000000000011011111001",
						 "100000000000011111111000",
						 "100000000000100011110111",
						 "100000000000100111110110",
						 "100000000000101011110101",
						 "100000000000101111110100",
						 "100000000000110011110011",
						 "100000000000110111110010",
						 "100000000000111011110001",
						 "100000000000000000000000",
						 "100000000000000011111111",
						 "100000000000000111111110",
						 "100000000000001011111101",
						 "100000000000001111111100",
						 "100000000000010011111011",
						 "100000000000010111111010",
						 "100000000000011011111001",
						 "100000000000011111111000",
						 "100000000000100011110111",
						 "100000000000100111110110",
						 "100000000000101011110101",
						 "100000000000101111110100",
						 "100000000000110011110011",
						 "100000000000110111110010",
						 "100000000000111011110001",
						 "100000000010100010111110",
						 "100000000010100110111101",
						 "100000000010101010111100",
						 "100000000010101110111011",
						 "100000000010110010111010",
						 "100000000010110110111001",
						 "100000000010111010111000",
						 "100000000010111110110111",
						 "100000000011000010110110",
						 "100000000011000110110101",
						 "100000000011001010110100",
						 "100000000011001110110011",
						 "100000000011010010110010",
						 "100000000011010110110001",
						 "100000000011011010110000",
						 "100000000011011110101111",
						 "100000000010100010111110",
						 "100000000010100110111101",
						 "100000000010101010111100",
						 "100000000010101110111011",
						 "100000000010110010111010",
						 "100000000010110110111001",
						 "100000000010111010111000",
						 "100000000010111110110111",
						 "100000000011000010110110",
						 "100000000011000110110101",
						 "100000000011001010110100",
						 "100000000011001110110011",
						 "100000000011010010110010",
						 "100000000011010110110001",
						 "100000000011011010110000",
						 "100000000011011110101111",
						 "100000000101000101111100",
						 "100000000101001001111011",
						 "100000000101001101111010",
						 "100000000101010001111001",
						 "100000000101010101111000",
						 "100000000101011001110111",
						 "100000000101011101110110",
						 "100000000101100001110101",
						 "100000000101100101110100",
						 "100000000101101001110011",
						 "100000000101101101110010",
						 "100000000101110001110001",
						 "100000000101110101110000",
						 "100000000101111001101111",
						 "100000000101111101101110",
						 "100000000110000001101101",
						 "100000000101000101111100",
						 "100000000101001001111011",
						 "100000000101001101111010",
						 "100000000101010001111001",
						 "100000000101010101111000",
						 "100000000101011001110111",
						 "100000000101011101110110",
						 "100000000101100001110101",
						 "100000000101100101110100",
						 "100000000101101001110011",
						 "100000000101101101110010",
						 "100000000101110001110001",
						 "100000000101110101110000",
						 "100000000101111001101111",
						 "100000000101111101101110",
						 "100000000110000001101101",
						 "100000000101000101111100",
						 "100000000101001001111011",
						 "100000000101001101111010",
						 "100000000101010001111001",
						 "100000000101010101111000",
						 "100000000101011001110111",
						 "100000000101011101110110",
						 "100000000101100001110101",
						 "100000000101100101110100",
						 "100000000101101001110011",
						 "100000000101101101110010",
						 "100000000101110001110001",
						 "100000000101110101110000",
						 "100000000101111001101111",
						 "100000000101111101101110",
						 "100000000110000001101101",
						 "100000000111101000111010",
						 "100000000111101100111001",
						 "100000000111110000111000",
						 "100000000111110100110111",
						 "100000000111111000110110",
						 "100000000111111100110101",
						 "100000001000000000110100",
						 "100000001000000100110011",
						 "100000001000001000110010",
						 "100000001000001100110001",
						 "100000001000010000110000",
						 "100000001000010100101111",
						 "100000001000011000101110",
						 "100000001000011100101101",
						 "100000001000100000101100",
						 "100000001000100100101011",
						 "100000000111101000111010",
						 "100000000111101100111001",
						 "100000000111110000111000",
						 "100000000111110100110111",
						 "100000000111111000110110",
						 "100000000111111100110101",
						 "100000001000000000110100",
						 "100000001000000100110011",
						 "100000001000001000110010",
						 "100000001000001100110001",
						 "100000001000010000110000",
						 "100000001000010100101111",
						 "100000001000011000101110",
						 "100000001000011100101101",
						 "100000001000100000101100",
						 "100000001000100100101011",
						 "100000001010001011111000",
						 "100000001010001111110111",
						 "100000001010010011110110",
						 "100000001010010111110101",
						 "100000001010011011110100",
						 "100000001010011111110011",
						 "100000001010100011110010",
						 "100000001010100111110001",
						 "100000001010101011110000",
						 "100000001010101111101111",
						 "100000001010110011101110",
						 "100000001010110111101101",
						 "100000001010111011101100",
						 "100000001010111111101011",
						 "100000001011000011101010",
						 "100000001011000111101001",
						 "100000001010001011111000",
						 "100000001010001111110111",
						 "100000001010010011110110",
						 "100000001010010111110101",
						 "100000001010011011110100",
						 "100000001010011111110011",
						 "100000001010100011110010",
						 "100000001010100111110001",
						 "100000001010101011110000",
						 "100000001010101111101111",
						 "100000001010110011101110",
						 "100000001010110111101101",
						 "100000001010111011101100",
						 "100000001010111111101011",
						 "100000001011000011101010",
						 "100000001011000111101001",
						 "100000001010001011111000",
						 "100000001010001111110111",
						 "100000001010010011110110",
						 "100000001010010111110101",
						 "100000001010011011110100",
						 "100000001010011111110011",
						 "100000001010100011110010",
						 "100000001010100111110001",
						 "100000001010101011110000",
						 "100000001010101111101111",
						 "100000001010110011101110",
						 "100000001010110111101101",
						 "100000001010111011101100",
						 "100000001010111111101011",
						 "100000001011000011101010",
						 "100000001011000111101001",
						 "100000001100101110110110",
						 "100000001100110010110101",
						 "100000001100110110110100",
						 "100000001100111010110011",
						 "100000001100111110110010",
						 "100000001101000010110001",
						 "100000001101000110110000",
						 "100000001101001010101111",
						 "100000001101001110101110",
						 "100000001101010010101101",
						 "100000001101010110101100",
						 "100000001101011010101011",
						 "100000001101011110101010",
						 "100000001101100010101001",
						 "100000001101100110101000",
						 "100000001101101010100111",
						 "100000001100101110110110",
						 "100000001100110010110101",
						 "100000001100110110110100",
						 "100000001100111010110011",
						 "100000001100111110110010",
						 "100000001101000010110001",
						 "100000001101000110110000",
						 "100000001101001010101111",
						 "100000001101001110101110",
						 "100000001101010010101101",
						 "100000001101010110101100",
						 "100000001101011010101011",
						 "100000001101011110101010",
						 "100000001101100010101001",
						 "100000001101100110101000",
						 "100000001101101010100111",
						 "100000001100101110110110",
						 "100000001100110010110101",
						 "100000001100110110110100",
						 "100000001100111010110011",
						 "100000001100111110110010",
						 "100000001101000010110001",
						 "100000001101000110110000",
						 "100000001101001010101111",
						 "100000001101001110101110",
						 "100000001101010010101101",
						 "100000001101010110101100",
						 "100000001101011010101011",
						 "100000001101011110101010",
						 "100000001101100010101001",
						 "100000001101100110101000",
						 "100000001101101010100111",
						 "100000001111010001110100",
						 "100000001111010101110011",
						 "100000001111011001110010",
						 "100000001111011101110001",
						 "100000001111100001110000",
						 "100000001111100101101111",
						 "100000001111101001101110",
						 "100000001111101101101101",
						 "100000001111110001101100",
						 "100000001111110101101011",
						 "100000001111111001101010",
						 "100000001111111101101001",
						 "100000010000000001101000",
						 "100000010000000101100111",
						 "100000010000001001100110",
						 "100000010000001101100101",
						 "100000001111010001110100",
						 "100000001111010101110011",
						 "100000001111011001110010",
						 "100000001111011101110001",
						 "100000001111100001110000",
						 "100000001111100101101111",
						 "100000001111101001101110",
						 "100000001111101101101101",
						 "100000001111110001101100",
						 "100000001111110101101011",
						 "100000001111111001101010",
						 "100000001111111101101001",
						 "100000010000000001101000",
						 "100000010000000101100111",
						 "100000010000001001100110",
						 "100000010000001101100101",
						 "100000010001110100110010",
						 "100000010001111000110001",
						 "100000010001111100110000",
						 "100000010010000000101111",
						 "100000010010000100101110",
						 "100000010010001000101101",
						 "100000010010001100101100",
						 "100000010010010000101011",
						 "100000010010010100101010",
						 "100000010010011000101001",
						 "100000010010011100101000",
						 "100000010010100000100111",
						 "100000010010100100100110",
						 "100000010010101000100101",
						 "100000010010101100100100",
						 "100000010010110000100011",
						 "100000010001110100110010",
						 "100000010001111000110001",
						 "100000010001111100110000",
						 "100000010010000000101111",
						 "100000010010000100101110",
						 "100000010010001000101101",
						 "100000010010001100101100",
						 "100000010010010000101011",
						 "100000010010010100101010",
						 "100000010010011000101001",
						 "100000010010011100101000",
						 "100000010010100000100111",
						 "100000010010100100100110",
						 "100000010010101000100101",
						 "100000010010101100100100",
						 "100000010010110000100011",
						 "100000010001110100110010",
						 "100000010001111000110001",
						 "100000010001111100110000",
						 "100000010010000000101111",
						 "100000010010000100101110",
						 "100000010010001000101101",
						 "100000010010001100101100",
						 "100000010010010000101011",
						 "100000010010010100101010",
						 "100000010010011000101001",
						 "100000010010011100101000",
						 "100000010010100000100111",
						 "100000010010100100100110",
						 "100000010010101000100101",
						 "100000010010101100100100",
						 "100000010010110000100011",
						 "100000010100010111110000",
						 "100000010100011011101111",
						 "100000010100011111101110",
						 "100000010100100011101101",
						 "100000010100100111101100",
						 "100000010100101011101011",
						 "100000010100101111101010",
						 "100000010100110011101001",
						 "100000010100110111101000",
						 "100000010100111011100111",
						 "100000010100111111100110",
						 "100000010101000011100101",
						 "100000010101000111100100",
						 "100000010101001011100011",
						 "100000010101001111100010",
						 "100000010101010011100001",
						 "100000010100010111110000",
						 "100000010100011011101111",
						 "100000010100011111101110",
						 "100000010100100011101101",
						 "100000010100100111101100",
						 "100000010100101011101011",
						 "100000010100101111101010",
						 "100000010100110011101001",
						 "100000010100110111101000",
						 "100000010100111011100111",
						 "100000010100111111100110",
						 "100000010101000011100101",
						 "100000010101000111100100",
						 "100000010101001011100011",
						 "100000010101001111100010",
						 "100000010101010011100001",
						 "100000010110111010101110",
						 "100000010110111110101101",
						 "100000010111000010101100",
						 "100000010111000110101011",
						 "100000010111001010101010",
						 "100000010111001110101001",
						 "100000010111010010101000",
						 "100000010111010110100111",
						 "100000010111011010100110",
						 "100000010111011110100101",
						 "100000010111100010100100",
						 "100000010111100110100011",
						 "100000010111101010100010",
						 "100000010111101110100001",
						 "100000010111110010100000",
						 "100000010111110110011111",
						 "100000010110111010101110",
						 "100000010110111110101101",
						 "100000010111000010101100",
						 "100000010111000110101011",
						 "100000010111001010101010",
						 "100000010111001110101001",
						 "100000010111010010101000",
						 "100000010111010110100111",
						 "100000010111011010100110",
						 "100000010111011110100101",
						 "100000010111100010100100",
						 "100000010111100110100011",
						 "100000010111101010100010",
						 "100000010111101110100001",
						 "100000010111110010100000",
						 "100000010111110110011111",
						 "100000010110111010101110",
						 "100000010110111110101101",
						 "100000010111000010101100",
						 "100000010111000110101011",
						 "100000010111001010101010",
						 "100000010111001110101001",
						 "100000010111010010101000",
						 "100000010111010110100111",
						 "100000010111011010100110",
						 "100000010111011110100101",
						 "100000010111100010100100",
						 "100000010111100110100011",
						 "100000010111101010100010",
						 "100000010111101110100001",
						 "100000010111110010100000",
						 "100000010111110110011111",
						 "100000011001011101101100",
						 "100000011001100001101011",
						 "100000011001100101101010",
						 "100000011001101001101001",
						 "100000011001101101101000",
						 "100000011001110001100111",
						 "100000011001110101100110",
						 "100000011001111001100101",
						 "100000011001111101100100",
						 "100000011010000001100011",
						 "100000011010000101100010",
						 "100000011010001001100001",
						 "100000011010001101100000",
						 "100000011010010001011111",
						 "100000011010010101011110",
						 "100000011010011001011101",
						 "100000011001011101101100",
						 "100000011001100001101011",
						 "100000011001100101101010",
						 "100000011001101001101001",
						 "100000011001101101101000",
						 "100000011001110001100111",
						 "100000011001110101100110",
						 "100000011001111001100101",
						 "100000011001111101100100",
						 "100000011010000001100011",
						 "100000011010000101100010",
						 "100000011010001001100001",
						 "100000011010001101100000",
						 "100000011010010001011111",
						 "100000011010010101011110",
						 "100000011010011001011101",
						 "100000011100000000101010",
						 "100000011100000100101001",
						 "100000011100001000101000",
						 "100000011100001100100111",
						 "100000011100010000100110",
						 "100000011100010100100101",
						 "100000011100011000100100",
						 "100000011100011100100011",
						 "100000011100100000100010",
						 "100000011100100100100001",
						 "100000011100101000100000",
						 "100000011100101100011111",
						 "100000011100110000011110",
						 "100000011100110100011101",
						 "100000011100111000011100",
						 "100000011100111100011011",
						 "100000011100000000101010",
						 "100000011100000100101001",
						 "100000011100001000101000",
						 "100000011100001100100111",
						 "100000011100010000100110",
						 "100000011100010100100101",
						 "100000011100011000100100",
						 "100000011100011100100011",
						 "100000011100100000100010",
						 "100000011100100100100001",
						 "100000011100101000100000",
						 "100000011100101100011111",
						 "100000011100110000011110",
						 "100000011100110100011101",
						 "100000011100111000011100",
						 "100000011100111100011011",
						 "100000011100000000101010",
						 "100000011100000100101001",
						 "100000011100001000101000",
						 "100000011100001100100111",
						 "100000011100010000100110",
						 "100000011100010100100101",
						 "100000011100011000100100",
						 "100000011100011100100011",
						 "100000011100100000100010",
						 "100000011100100100100001",
						 "100000011100101000100000",
						 "100000011100101100011111",
						 "100000011100110000011110",
						 "100000011100110100011101",
						 "100000011100111000011100",
						 "100000011100111100011011",
						 "100000011110100011101000",
						 "100000011110100111100111",
						 "100000011110101011100110",
						 "100000011110101111100101",
						 "100000011110110011100100",
						 "100000011110110111100011",
						 "100000011110111011100010",
						 "100000011110111111100001",
						 "100000011111000011100000",
						 "100000011111000111011111",
						 "100000011111001011011110",
						 "100000011111001111011101",
						 "100000011111010011011100",
						 "100000011111010111011011",
						 "100000011111011011011010",
						 "100000011111011111011001",
						 "100000011110100011101000",
						 "100000011110100111100111",
						 "100000011110101011100110",
						 "100000011110101111100101",
						 "100000011110110011100100",
						 "100000011110110111100011",
						 "100000011110111011100010",
						 "100000011110111111100001",
						 "100000011111000011100000",
						 "100000011111000111011111",
						 "100000011111001011011110",
						 "100000011111001111011101",
						 "100000011111010011011100",
						 "100000011111010111011011",
						 "100000011111011011011010",
						 "100000011111011111011001",
						 "100000100001000110100110",
						 "100000100001001010100101",
						 "100000100001001110100100",
						 "100000100001010010100011",
						 "100000100001010110100010",
						 "100000100001011010100001",
						 "100000100001011110100000",
						 "100000100001100010011111",
						 "100000100001100110011110",
						 "100000100001101010011101",
						 "100000100001101110011100",
						 "100000100001110010011011",
						 "100000100001110110011010",
						 "100000100001111010011001",
						 "100000100001111110011000",
						 "100000100010000010010111",
						 "100000100001000110100110",
						 "100000100001001010100101",
						 "100000100001001110100100",
						 "100000100001010010100011",
						 "100000100001010110100010",
						 "100000100001011010100001",
						 "100000100001011110100000",
						 "100000100001100010011111",
						 "100000100001100110011110",
						 "100000100001101010011101",
						 "100000100001101110011100",
						 "100000100001110010011011",
						 "100000100001110110011010",
						 "100000100001111010011001",
						 "100000100001111110011000",
						 "100000100010000010010111",
						 "100000100001000110100110",
						 "100000100001001010100101",
						 "100000100001001110100100",
						 "100000100001010010100011",
						 "100000100001010110100010",
						 "100000100001011010100001",
						 "100000100001011110100000",
						 "100000100001100010011111",
						 "100000100001100110011110",
						 "100000100001101010011101",
						 "100000100001101110011100",
						 "100000100001110010011011",
						 "100000100001110110011010",
						 "100000100001111010011001",
						 "100000100001111110011000",
						 "100000100010000010010111",
						 "100000100011101001100100",
						 "100000100011101101100011",
						 "100000100011110001100010",
						 "100000100011110101100001",
						 "100000100011111001100000",
						 "100000100011111101011111",
						 "100000100100000001011110",
						 "100000100100000101011101",
						 "100000100100001001011100",
						 "100000100100001101011011",
						 "100000100100010001011010",
						 "100000100100010101011001",
						 "100000100100011001011000",
						 "100000100100011101010111",
						 "100000100100100001010110",
						 "100000100100100101010101",
						 "100000100011101001100100",
						 "100000100011101101100011",
						 "100000100011110001100010",
						 "100000100011110101100001",
						 "100000100011111001100000",
						 "100000100011111101011111",
						 "100000100100000001011110",
						 "100000100100000101011101",
						 "100000100100001001011100",
						 "100000100100001101011011",
						 "100000100100010001011010",
						 "100000100100010101011001",
						 "100000100100011001011000",
						 "100000100100011101010111",
						 "100000100100100001010110",
						 "100000100100100101010101",
						 "100000100011101001100100",
						 "100000100011101101100011",
						 "100000100011110001100010",
						 "100000100011110101100001",
						 "100000100011111001100000",
						 "100000100011111101011111",
						 "100000100100000001011110",
						 "100000100100000101011101",
						 "100000100100001001011100",
						 "100000100100001101011011",
						 "100000100100010001011010",
						 "100000100100010101011001",
						 "100000100100011001011000",
						 "100000100100011101010111",
						 "100000100100100001010110",
						 "100000100100100101010101",
						 "100000100110001100100010",
						 "100000100110010000100001",
						 "100000100110010100100000",
						 "100000100110011000011111",
						 "100000100110011100011110",
						 "100000100110100000011101",
						 "100000100110100100011100",
						 "100000100110101000011011",
						 "100000100110101100011010",
						 "100000100110110000011001",
						 "100000100110110100011000",
						 "100000100110111000010111",
						 "100000100110111100010110",
						 "100000100111000000010101",
						 "100000100111000100010100",
						 "100000100111001000010011",
						 "100000100110001100100010",
						 "100000100110010000100001",
						 "100000100110010100100000",
						 "100000100110011000011111",
						 "100000100110011100011110",
						 "100000100110100000011101",
						 "100000100110100100011100",
						 "100000100110101000011011",
						 "100000100110101100011010",
						 "100000100110110000011001",
						 "100000100110110100011000",
						 "100000100110111000010111",
						 "100000100110111100010110",
						 "100000100111000000010101",
						 "100000100111000100010100",
						 "100000100111001000010011",
						 "100000101000101111100000",
						 "100000101000110011011111",
						 "100000101000110111011110",
						 "100000101000111011011101",
						 "100000101000111111011100",
						 "100000101001000011011011",
						 "100000101001000111011010",
						 "100000101001001011011001",
						 "100000101001001111011000",
						 "100000101001010011010111",
						 "100000101001010111010110",
						 "100000101001011011010101",
						 "100000101001011111010100",
						 "100000101001100011010011",
						 "100000101001100111010010",
						 "100000101001101011010001",
						 "100000101000101111100000",
						 "100000101000110011011110",
						 "100000101000110111011100",
						 "100000101000111011011010",
						 "100000101000111111011000",
						 "100000101001000011010110",
						 "100000101001000111010100",
						 "100000101001001011010010",
						 "100000101001001111010000",
						 "100000101001010011001110",
						 "100000101001010111001100",
						 "100000101001011011001010",
						 "100000101001011111001000",
						 "100000101001100011000110",
						 "100000101001100111000100",
						 "100000101001101011000010",
						 "100000101000101111100000",
						 "100000101000110011011110",
						 "100000101000110111011100",
						 "100000101000111011011010",
						 "100000101000111111011000",
						 "100000101001000011010110",
						 "100000101001000111010100",
						 "100000101001001011010010",
						 "100000101001001111010000",
						 "100000101001010011001110",
						 "100000101001010111001100",
						 "100000101001011011001010",
						 "100000101001011111001000",
						 "100000101001100011000110",
						 "100000101001100111000100",
						 "100000101001101011000010",
						 "100000101011010010011110",
						 "100000101011010110011100",
						 "100000101011011010011010",
						 "100000101011011110011000",
						 "100000101011100010010110",
						 "100000101011100110010100",
						 "100000101011101010010010",
						 "100000101011101110010000",
						 "100000101011110010001110",
						 "100000101011110110001100",
						 "100000101011111010001010",
						 "100000101011111110001000",
						 "100000101100000010000110",
						 "100000101100000110000100",
						 "100000101100001010000010",
						 "100000101100001110000000",
						 "100000101011010010011110",
						 "100000101011010110011100",
						 "100000101011011010011010",
						 "100000101011011110011000",
						 "100000101011100010010110",
						 "100000101011100110010100",
						 "100000101011101010010010",
						 "100000101011101110010000",
						 "100000101011110010001110",
						 "100000101011110110001100",
						 "100000101011111010001010",
						 "100000101011111110001000",
						 "100000101100000010000110",
						 "100000101100000110000100",
						 "100000101100001010000010",
						 "100000101100001110000000",
						 "100000101101110101011100",
						 "100000101101111001011010",
						 "100000101101111101011000",
						 "100000101110000001010110",
						 "100000101110000101010100",
						 "100000101110001001010010",
						 "100000101110001101010000",
						 "100000101110010001001110",
						 "100000101110010101001100",
						 "100000101110011001001010",
						 "100000101110011101001000",
						 "100000101110100001000110",
						 "100000101110100101000100",
						 "100000101110101001000010",
						 "100000101110101101000000",
						 "100000101110110000111110",
						 "100000101101110101011100",
						 "100000101101111001011010",
						 "100000101101111101011000",
						 "100000101110000001010110",
						 "100000101110000101010100",
						 "100000101110001001010010",
						 "100000101110001101010000",
						 "100000101110010001001110",
						 "100000101110010101001100",
						 "100000101110011001001010",
						 "100000101110011101001000",
						 "100000101110100001000110",
						 "100000101110100101000100",
						 "100000101110101001000010",
						 "100000101110101101000000",
						 "100000101110110000111110",
						 "100000101101110101011100",
						 "100000101101111001011010",
						 "100000101101111101011000",
						 "100000101110000001010110",
						 "100000101110000101010100",
						 "100000101110001001010010",
						 "100000101110001101010000",
						 "100000101110010001001110",
						 "100000101110010101001100",
						 "100000101110011001001010",
						 "100000101110011101001000",
						 "100000101110100001000110",
						 "100000101110100101000100",
						 "100000101110101001000010",
						 "100000101110101101000000",
						 "100000101110110000111110",
						 "100000110000011000011010",
						 "100000110000011100011000",
						 "100000110000100000010110",
						 "100000110000100100010100",
						 "100000110000101000010010",
						 "100000110000101100010000",
						 "100000110000110000001110",
						 "100000110000110100001100",
						 "100000110000111000001010",
						 "100000110000111100001000",
						 "100000110001000000000110",
						 "100000110001000100000100",
						 "100000110001001000000010",
						 "100000110001001100000000",
						 "100000110001001111111110",
						 "100000110001010011111100",
						 "100000110000011000011010",
						 "100000110000011100011000",
						 "100000110000100000010110",
						 "100000110000100100010100",
						 "100000110000101000010010",
						 "100000110000101100010000",
						 "100000110000110000001110",
						 "100000110000110100001100",
						 "100000110000111000001010",
						 "100000110000111100001000",
						 "100000110001000000000110",
						 "100000110001000100000100",
						 "100000110001001000000010",
						 "100000110001001100000000",
						 "100000110001001111111110",
						 "100000110001010011111100",
						 "100000110010111011011000",
						 "100000110010111111010110",
						 "100000110011000011010100",
						 "100000110011000111010010",
						 "100000110011001011010000",
						 "100000110011001111001110",
						 "100000110011010011001100",
						 "100000110011010111001010",
						 "100000110011011011001000",
						 "100000110011011111000110",
						 "100000110011100011000100",
						 "100000110011100111000010",
						 "100000110011101011000000",
						 "100000110011101110111110",
						 "100000110011110010111100",
						 "100000110011110110111010",
						 "100000110010111011011000",
						 "100000110010111111010110",
						 "100000110011000011010100",
						 "100000110011000111010010",
						 "100000110011001011010000",
						 "100000110011001111001110",
						 "100000110011010011001100",
						 "100000110011010111001010",
						 "100000110011011011001000",
						 "100000110011011111000110",
						 "100000110011100011000100",
						 "100000110011100111000010",
						 "100000110011101011000000",
						 "100000110011101110111110",
						 "100000110011110010111100",
						 "100000110011110110111010",
						 "100000110010111011011000",
						 "100000110010111111010110",
						 "100000110011000011010100",
						 "100000110011000111010010",
						 "100000110011001011010000",
						 "100000110011001111001110",
						 "100000110011010011001100",
						 "100000110011010111001010",
						 "100000110011011011001000",
						 "100000110011011111000110",
						 "100000110011100011000100",
						 "100000110011100111000010",
						 "100000110011101011000000",
						 "100000110011101110111110",
						 "100000110011110010111100",
						 "100000110011110110111010",
						 "100000110101011110010110",
						 "100000110101100010010100",
						 "100000110101100110010010",
						 "100000110101101010010000",
						 "100000110101101110001110",
						 "100000110101110010001100",
						 "100000110101110110001010",
						 "100000110101111010001000",
						 "100000110101111110000110",
						 "100000110110000010000100",
						 "100000110110000110000010",
						 "100000110110001010000000",
						 "100000110110001101111110",
						 "100000110110010001111100",
						 "100000110110010101111010",
						 "100000110110011001111000",
						 "100000110101011110010110",
						 "100000110101100010010100",
						 "100000110101100110010010",
						 "100000110101101010010000",
						 "100000110101101110001110",
						 "100000110101110010001100",
						 "100000110101110110001010",
						 "100000110101111010001000",
						 "100000110101111110000110",
						 "100000110110000010000100",
						 "100000110110000110000010",
						 "100000110110001010000000",
						 "100000110110001101111110",
						 "100000110110010001111100",
						 "100000110110010101111010",
						 "100000110110011001111000",
						 "100000110101011110010110",
						 "100000110101100010010100",
						 "100000110101100110010010",
						 "100000110101101010010000",
						 "100000110101101110001110",
						 "100000110101110010001100",
						 "100000110101110110001010",
						 "100000110101111010001000",
						 "100000110101111110000110",
						 "100000110110000010000100",
						 "100000110110000110000010",
						 "100000110110001010000000",
						 "100000110110001101111110",
						 "100000110110010001111100",
						 "100000110110010101111010",
						 "100000110110011001111000",
						 "100000111000000001010100",
						 "100000111000000101010010",
						 "100000111000001001010000",
						 "100000111000001101001110",
						 "100000111000010001001100",
						 "100000111000010101001010",
						 "100000111000011001001000",
						 "100000111000011101000110",
						 "100000111000100001000100",
						 "100000111000100101000010",
						 "100000111000101001000000",
						 "100000111000101100111110",
						 "100000111000110000111100",
						 "100000111000110100111010",
						 "100000111000111000111000",
						 "100000111000111100110110",
						 "100000111000000001010100",
						 "100000111000000101010010",
						 "100000111000001001010000",
						 "100000111000001101001110",
						 "100000111000010001001100",
						 "100000111000010101001010",
						 "100000111000011001001000",
						 "100000111000011101000110",
						 "100000111000100001000100",
						 "100000111000100101000010",
						 "100000111000101001000000",
						 "100000111000101100111110",
						 "100000111000110000111100",
						 "100000111000110100111010",
						 "100000111000111000111000",
						 "100000111000111100110110",
						 "100000111010100100010010",
						 "100000111010101000010000",
						 "100000111010101100001110",
						 "100000111010110000001100",
						 "100000111010110100001010",
						 "100000111010111000001000",
						 "100000111010111100000110",
						 "100000111011000000000100",
						 "100000111011000100000010",
						 "100000111011001000000000",
						 "100000111011001011111110",
						 "100000111011001111111100",
						 "100000111011010011111010",
						 "100000111011010111111000",
						 "100000111011011011110110",
						 "100000111011011111110100",
						 "100000111010100100010010",
						 "100000111010101000010000",
						 "100000111010101100001110",
						 "100000111010110000001100",
						 "100000111010110100001010",
						 "100000111010111000001000",
						 "100000111010111100000110",
						 "100000111011000000000100",
						 "100000111011000100000010",
						 "100000111011001000000000",
						 "100000111011001011111110",
						 "100000111011001111111100",
						 "100000111011010011111010",
						 "100000111011010111111000",
						 "100000111011011011110110",
						 "100000111011011111110100",
						 "100000111010100100010010",
						 "100000111010101000010000",
						 "100000111010101100001110",
						 "100000111010110000001100",
						 "100000111010110100001010",
						 "100000111010111000001000",
						 "100000111010111100000110",
						 "100000111011000000000100",
						 "100000111011000100000010",
						 "100000111011001000000000",
						 "100000111011001011111110",
						 "100000111011001111111100",
						 "100000111011010011111010",
						 "100000111011010111111000",
						 "100000111011011011110110",
						 "100000111011011111110100",
						 "100000111101000111010000",
						 "100000111101001011001110",
						 "100000111101001111001100",
						 "100000111101010011001010",
						 "100000111101010111001000",
						 "100000111101011011000110",
						 "100000111101011111000100",
						 "100000111101100011000010",
						 "100000111101100111000000",
						 "100000111101101010111110",
						 "100000111101101110111100",
						 "100000111101110010111010",
						 "100000111101110110111000",
						 "100000111101111010110110",
						 "100000111101111110110100",
						 "100000111110000010110010",
						 "100000111101000111010000",
						 "100000111101001011001110",
						 "100000111101001111001100",
						 "100000111101010011001010",
						 "100000111101010111001000",
						 "100000111101011011000110",
						 "100000111101011111000100",
						 "100000111101100011000010",
						 "100000111101100111000000",
						 "100000111101101010111110",
						 "100000111101101110111100",
						 "100000111101110010111010",
						 "100000111101110110111000",
						 "100000111101111010110110",
						 "100000111101111110110100",
						 "100000111110000010110010",
						 "100000111111101010001110",
						 "100000111111101110001100",
						 "100000111111110010001010",
						 "100000111111110110001000",
						 "100000111111111010000110",
						 "100000111111111110000100",
						 "100001000000000010000010",
						 "100001000000000110000000",
						 "100001000000001001111110",
						 "100001000000001101111100",
						 "100001000000010001111010",
						 "100001000000010101111000",
						 "100001000000011001110110",
						 "100001000000011101110100",
						 "100001000000100001110010",
						 "100001000000100101110000",
						 "100000111111101010001110",
						 "100000111111101110001100",
						 "100000111111110010001010",
						 "100000111111110110001000",
						 "100000111111111010000110",
						 "100000111111111110000100",
						 "100001000000000010000010",
						 "100001000000000110000000",
						 "100001000000001001111110",
						 "100001000000001101111100",
						 "100001000000010001111010",
						 "100001000000010101111000",
						 "100001000000011001110110",
						 "100001000000011101110100",
						 "100001000000100001110010",
						 "100001000000100101110000",
						 "100000111111101010001110",
						 "100000111111101110001100",
						 "100000111111110010001010",
						 "100000111111110110001000",
						 "100000111111111010000110",
						 "100000111111111110000100",
						 "100001000000000010000010",
						 "100001000000000110000000",
						 "100001000000001001111110",
						 "100001000000001101111100",
						 "100001000000010001111010",
						 "100001000000010101111000",
						 "100001000000011001110110",
						 "100001000000011101110100",
						 "100001000000100001110010",
						 "100001000000100101110000",
						 "100001000010001101001100",
						 "100001000010010001001010",
						 "100001000010010101001000",
						 "100001000010011001000110",
						 "100001000010011101000100",
						 "100001000010100001000010",
						 "100001000010100101000000",
						 "100001000010101000111110",
						 "100001000010101100111100",
						 "100001000010110000111010",
						 "100001000010110100111000",
						 "100001000010111000110110",
						 "100001000010111100110100",
						 "100001000011000000110010",
						 "100001000011000100110000",
						 "100001000011001000101110",
						 "100001000010001101001100",
						 "100001000010010001001010",
						 "100001000010010101001000",
						 "100001000010011001000110",
						 "100001000010011101000100",
						 "100001000010100001000010",
						 "100001000010100101000000",
						 "100001000010101000111110",
						 "100001000010101100111100",
						 "100001000010110000111010",
						 "100001000010110100111000",
						 "100001000010111000110110",
						 "100001000010111100110100",
						 "100001000011000000110010",
						 "100001000011000100110000",
						 "100001000011001000101110",
						 "100001000100110000001010",
						 "100001000100110100001000",
						 "100001000100111000000110",
						 "100001000100111100000100",
						 "100001000101000000000010",
						 "100001000101000100000000",
						 "100001000101000111111110",
						 "100001000101001011111100",
						 "100001000101001111111010",
						 "100001000101010011111000",
						 "100001000101010111110110",
						 "100001000101011011110100",
						 "100001000101011111110010",
						 "100001000101100011110000",
						 "100001000101100111101110",
						 "100001000101101011101100",
						 "100001000100110000001010",
						 "100001000100110100001000",
						 "100001000100111000000110",
						 "100001000100111100000100",
						 "100001000101000000000010",
						 "100001000101000100000000",
						 "100001000101000111111110",
						 "100001000101001011111100",
						 "100001000101001111111010",
						 "100001000101010011111000",
						 "100001000101010111110110",
						 "100001000101011011110100",
						 "100001000101011111110010",
						 "100001000101100011110000",
						 "100001000101100111101110",
						 "100001000101101011101100",
						 "100001000100110000001010",
						 "100001000100110100001000",
						 "100001000100111000000110",
						 "100001000100111100000100",
						 "100001000101000000000010",
						 "100001000101000100000000",
						 "100001000101000111111110",
						 "100001000101001011111100",
						 "100001000101001111111010",
						 "100001000101010011111000",
						 "100001000101010111110110",
						 "100001000101011011110100",
						 "100001000101011111110010",
						 "100001000101100011110000",
						 "100001000101100111101110",
						 "100001000101101011101100",
						 "100001000111010011001000",
						 "100001000111010111000101",
						 "100001000111011011000010",
						 "100001000111011110111111",
						 "100001000111100010111100",
						 "100001000111100110111001",
						 "100001000111101010110110",
						 "100001000111101110110011",
						 "100001000111110010110000",
						 "100001000111110110101101",
						 "100001000111111010101010",
						 "100001000111111110100111",
						 "100001001000000010100100",
						 "100001001000000110100001",
						 "100001001000001010011110",
						 "100001001000001110011011",
						 "100001000111010011001000",
						 "100001000111010111000101",
						 "100001000111011011000010",
						 "100001000111011110111111",
						 "100001000111100010111100",
						 "100001000111100110111001",
						 "100001000111101010110110",
						 "100001000111101110110011",
						 "100001000111110010110000",
						 "100001000111110110101101",
						 "100001000111111010101010",
						 "100001000111111110100111",
						 "100001001000000010100100",
						 "100001001000000110100001",
						 "100001001000001010011110",
						 "100001001000001110011011",
						 "100001000111010011001000",
						 "100001000111010111000101",
						 "100001000111011011000010",
						 "100001000111011110111111",
						 "100001000111100010111100",
						 "100001000111100110111001",
						 "100001000111101010110110",
						 "100001000111101110110011",
						 "100001000111110010110000",
						 "100001000111110110101101",
						 "100001000111111010101010",
						 "100001000111111110100111",
						 "100001001000000010100100",
						 "100001001000000110100001",
						 "100001001000001010011110",
						 "100001001000001110011011",
						 "100001001001110110000110",
						 "100001001001111010000011",
						 "100001001001111110000000",
						 "100001001010000001111101",
						 "100001001010000101111010",
						 "100001001010001001110111",
						 "100001001010001101110100",
						 "100001001010010001110001",
						 "100001001010010101101110",
						 "100001001010011001101011",
						 "100001001010011101101000",
						 "100001001010100001100101",
						 "100001001010100101100010",
						 "100001001010101001011111",
						 "100001001010101101011100",
						 "100001001010110001011001",
						 "100001001001110110000110",
						 "100001001001111010000011",
						 "100001001001111110000000",
						 "100001001010000001111101",
						 "100001001010000101111010",
						 "100001001010001001110111",
						 "100001001010001101110100",
						 "100001001010010001110001",
						 "100001001010010101101110",
						 "100001001010011001101011",
						 "100001001010011101101000",
						 "100001001010100001100101",
						 "100001001010100101100010",
						 "100001001010101001011111",
						 "100001001010101101011100",
						 "100001001010110001011001",
						 "100001001100011001000100",
						 "100001001100011101000001",
						 "100001001100100000111110",
						 "100001001100100100111011",
						 "100001001100101000111000",
						 "100001001100101100110101",
						 "100001001100110000110010",
						 "100001001100110100101111",
						 "100001001100111000101100",
						 "100001001100111100101001",
						 "100001001101000000100110",
						 "100001001101000100100011",
						 "100001001101001000100000",
						 "100001001101001100011101",
						 "100001001101010000011010",
						 "100001001101010100010111",
						 "100001001100011001000100",
						 "100001001100011101000001",
						 "100001001100100000111110",
						 "100001001100100100111011",
						 "100001001100101000111000",
						 "100001001100101100110101",
						 "100001001100110000110010",
						 "100001001100110100101111",
						 "100001001100111000101100",
						 "100001001100111100101001",
						 "100001001101000000100110",
						 "100001001101000100100011",
						 "100001001101001000100000",
						 "100001001101001100011101",
						 "100001001101010000011010",
						 "100001001101010100010111",
						 "100001001100011001000100",
						 "100001001100011101000001",
						 "100001001100100000111110",
						 "100001001100100100111011",
						 "100001001100101000111000",
						 "100001001100101100110101",
						 "100001001100110000110010",
						 "100001001100110100101111",
						 "100001001100111000101100",
						 "100001001100111100101001",
						 "100001001101000000100110",
						 "100001001101000100100011",
						 "100001001101001000100000",
						 "100001001101001100011101",
						 "100001001101010000011010",
						 "100001001101010100010111",
						 "100001001110111100000010",
						 "100001001110111111111111",
						 "100001001111000011111100",
						 "100001001111000111111001",
						 "100001001111001011110110",
						 "100001001111001111110011",
						 "100001001111010011110000",
						 "100001001111010111101101",
						 "100001001111011011101010",
						 "100001001111011111100111",
						 "100001001111100011100100",
						 "100001001111100111100001",
						 "100001001111101011011110",
						 "100001001111101111011011",
						 "100001001111110011011000",
						 "100001001111110111010101",
						 "100001001110111100000010",
						 "100001001110111111111111",
						 "100001001111000011111100",
						 "100001001111000111111001",
						 "100001001111001011110110",
						 "100001001111001111110011",
						 "100001001111010011110000",
						 "100001001111010111101101",
						 "100001001111011011101010",
						 "100001001111011111100111",
						 "100001001111100011100100",
						 "100001001111100111100001",
						 "100001001111101011011110",
						 "100001001111101111011011",
						 "100001001111110011011000",
						 "100001001111110111010101",
						 "100001010001011111000000",
						 "100001010001100010111101",
						 "100001010001100110111010",
						 "100001010001101010110111",
						 "100001010001101110110100",
						 "100001010001110010110001",
						 "100001010001110110101110",
						 "100001010001111010101011",
						 "100001010001111110101000",
						 "100001010010000010100101",
						 "100001010010000110100010",
						 "100001010010001010011111",
						 "100001010010001110011100",
						 "100001010010010010011001",
						 "100001010010010110010110",
						 "100001010010011010010011",
						 "100001010001011111000000",
						 "100001010001100010111101",
						 "100001010001100110111010",
						 "100001010001101010110111",
						 "100001010001101110110100",
						 "100001010001110010110001",
						 "100001010001110110101110",
						 "100001010001111010101011",
						 "100001010001111110101000",
						 "100001010010000010100101",
						 "100001010010000110100010",
						 "100001010010001010011111",
						 "100001010010001110011100",
						 "100001010010010010011001",
						 "100001010010010110010110",
						 "100001010010011010010011",
						 "100001010001011111000000",
						 "100001010001100010111101",
						 "100001010001100110111010",
						 "100001010001101010110111",
						 "100001010001101110110100",
						 "100001010001110010110001",
						 "100001010001110110101110",
						 "100001010001111010101011",
						 "100001010001111110101000",
						 "100001010010000010100101",
						 "100001010010000110100010",
						 "100001010010001010011111",
						 "100001010010001110011100",
						 "100001010010010010011001",
						 "100001010010010110010110",
						 "100001010010011010010011",
						 "100001010100000001111110",
						 "100001010100000101111011",
						 "100001010100001001111000",
						 "100001010100001101110101",
						 "100001010100010001110010",
						 "100001010100010101101111",
						 "100001010100011001101100",
						 "100001010100011101101001",
						 "100001010100100001100110",
						 "100001010100100101100011",
						 "100001010100101001100000",
						 "100001010100101101011101",
						 "100001010100110001011010",
						 "100001010100110101010111",
						 "100001010100111001010100",
						 "100001010100111101010001",
						 "100001010100000001111110",
						 "100001010100000101111011",
						 "100001010100001001111000",
						 "100001010100001101110101",
						 "100001010100010001110010",
						 "100001010100010101101111",
						 "100001010100011001101100",
						 "100001010100011101101001",
						 "100001010100100001100110",
						 "100001010100100101100011",
						 "100001010100101001100000",
						 "100001010100101101011101",
						 "100001010100110001011010",
						 "100001010100110101010111",
						 "100001010100111001010100",
						 "100001010100111101010001",
						 "100001010110100100111100",
						 "100001010110101000111001",
						 "100001010110101100110110",
						 "100001010110110000110011",
						 "100001010110110100110000",
						 "100001010110111000101101",
						 "100001010110111100101010",
						 "100001010111000000100111",
						 "100001010111000100100100",
						 "100001010111001000100001",
						 "100001010111001100011110",
						 "100001010111010000011011",
						 "100001010111010100011000",
						 "100001010111011000010101",
						 "100001010111011100010010",
						 "100001010111100000001111",
						 "100001010110100100111100",
						 "100001010110101000111001",
						 "100001010110101100110110",
						 "100001010110110000110011",
						 "100001010110110100110000",
						 "100001010110111000101101",
						 "100001010110111100101010",
						 "100001010111000000100111",
						 "100001010111000100100100",
						 "100001010111001000100001",
						 "100001010111001100011110",
						 "100001010111010000011011",
						 "100001010111010100011000",
						 "100001010111011000010101",
						 "100001010111011100010010",
						 "100001010111100000001111",
						 "100001010110100100111100",
						 "100001010110101000111001",
						 "100001010110101100110110",
						 "100001010110110000110011",
						 "100001010110110100110000",
						 "100001010110111000101101",
						 "100001010110111100101010",
						 "100001010111000000100111",
						 "100001010111000100100100",
						 "100001010111001000100001",
						 "100001010111001100011110",
						 "100001010111010000011011",
						 "100001010111010100011000",
						 "100001010111011000010101",
						 "100001010111011100010010",
						 "100001010111100000001111",
						 "100001011001000111111010",
						 "100001011001001011110111",
						 "100001011001001111110100",
						 "100001011001010011110001",
						 "100001011001010111101110",
						 "100001011001011011101011",
						 "100001011001011111101000",
						 "100001011001100011100101",
						 "100001011001100111100010",
						 "100001011001101011011111",
						 "100001011001101111011100",
						 "100001011001110011011001",
						 "100001011001110111010110",
						 "100001011001111011010011",
						 "100001011001111111010000",
						 "100001011010000011001101",
						 "100001011001000111111010",
						 "100001011001001011110111",
						 "100001011001001111110100",
						 "100001011001010011110001",
						 "100001011001010111101110",
						 "100001011001011011101011",
						 "100001011001011111101000",
						 "100001011001100011100101",
						 "100001011001100111100010",
						 "100001011001101011011111",
						 "100001011001101111011100",
						 "100001011001110011011001",
						 "100001011001110111010110",
						 "100001011001111011010011",
						 "100001011001111111010000",
						 "100001011010000011001101",
						 "100001011001000111111010",
						 "100001011001001011110110",
						 "100001011001001111110010",
						 "100001011001010011101110",
						 "100001011001010111101010",
						 "100001011001011011100110",
						 "100001011001011111100010",
						 "100001011001100011011110",
						 "100001011001100111011010",
						 "100001011001101011010110",
						 "100001011001101111010010",
						 "100001011001110011001110",
						 "100001011001110111001010",
						 "100001011001111011000110",
						 "100001011001111111000010",
						 "100001011010000010111110",
						 "100001011011101010111000",
						 "100001011011101110110100",
						 "100001011011110010110000",
						 "100001011011110110101100",
						 "100001011011111010101000",
						 "100001011011111110100100",
						 "100001011100000010100000",
						 "100001011100000110011100",
						 "100001011100001010011000",
						 "100001011100001110010100",
						 "100001011100010010010000",
						 "100001011100010110001100",
						 "100001011100011010001000",
						 "100001011100011110000100",
						 "100001011100100010000000",
						 "100001011100100101111100",
						 "100001011011101010111000",
						 "100001011011101110110100",
						 "100001011011110010110000",
						 "100001011011110110101100",
						 "100001011011111010101000",
						 "100001011011111110100100",
						 "100001011100000010100000",
						 "100001011100000110011100",
						 "100001011100001010011000",
						 "100001011100001110010100",
						 "100001011100010010010000",
						 "100001011100010110001100",
						 "100001011100011010001000",
						 "100001011100011110000100",
						 "100001011100100010000000",
						 "100001011100100101111100",
						 "100001011110001101110110",
						 "100001011110010001110010",
						 "100001011110010101101110",
						 "100001011110011001101010",
						 "100001011110011101100110",
						 "100001011110100001100010",
						 "100001011110100101011110",
						 "100001011110101001011010",
						 "100001011110101101010110",
						 "100001011110110001010010",
						 "100001011110110101001110",
						 "100001011110111001001010",
						 "100001011110111101000110",
						 "100001011111000001000010",
						 "100001011111000100111110",
						 "100001011111001000111010",
						 "100001011110001101110110",
						 "100001011110010001110010",
						 "100001011110010101101110",
						 "100001011110011001101010",
						 "100001011110011101100110",
						 "100001011110100001100010",
						 "100001011110100101011110",
						 "100001011110101001011010",
						 "100001011110101101010110",
						 "100001011110110001010010",
						 "100001011110110101001110",
						 "100001011110111001001010",
						 "100001011110111101000110",
						 "100001011111000001000010",
						 "100001011111000100111110",
						 "100001011111001000111010",
						 "100001011110001101110110",
						 "100001011110010001110010",
						 "100001011110010101101110",
						 "100001011110011001101010",
						 "100001011110011101100110",
						 "100001011110100001100010",
						 "100001011110100101011110",
						 "100001011110101001011010",
						 "100001011110101101010110",
						 "100001011110110001010010",
						 "100001011110110101001110",
						 "100001011110111001001010",
						 "100001011110111101000110",
						 "100001011111000001000010",
						 "100001011111000100111110",
						 "100001011111001000111010",
						 "100001100000110000110100",
						 "100001100000110100110000",
						 "100001100000111000101100",
						 "100001100000111100101000",
						 "100001100001000000100100",
						 "100001100001000100100000",
						 "100001100001001000011100",
						 "100001100001001100011000",
						 "100001100001010000010100",
						 "100001100001010100010000",
						 "100001100001011000001100",
						 "100001100001011100001000",
						 "100001100001100000000100",
						 "100001100001100100000000",
						 "100001100001100111111100",
						 "100001100001101011111000",
						 "100001100000110000110100",
						 "100001100000110100110000",
						 "100001100000111000101100",
						 "100001100000111100101000",
						 "100001100001000000100100",
						 "100001100001000100100000",
						 "100001100001001000011100",
						 "100001100001001100011000",
						 "100001100001010000010100",
						 "100001100001010100010000",
						 "100001100001011000001100",
						 "100001100001011100001000",
						 "100001100001100000000100",
						 "100001100001100100000000",
						 "100001100001100111111100",
						 "100001100001101011111000",
						 "100001100011010011110010",
						 "100001100011010111101110",
						 "100001100011011011101010",
						 "100001100011011111100110",
						 "100001100011100011100010",
						 "100001100011100111011110",
						 "100001100011101011011010",
						 "100001100011101111010110",
						 "100001100011110011010010",
						 "100001100011110111001110",
						 "100001100011111011001010",
						 "100001100011111111000110",
						 "100001100100000011000010",
						 "100001100100000110111110",
						 "100001100100001010111010",
						 "100001100100001110110110",
						 "100001100011010011110010",
						 "100001100011010111101110",
						 "100001100011011011101010",
						 "100001100011011111100110",
						 "100001100011100011100010",
						 "100001100011100111011110",
						 "100001100011101011011010",
						 "100001100011101111010110",
						 "100001100011110011010010",
						 "100001100011110111001110",
						 "100001100011111011001010",
						 "100001100011111111000110",
						 "100001100100000011000010",
						 "100001100100000110111110",
						 "100001100100001010111010",
						 "100001100100001110110110",
						 "100001100011010011110010",
						 "100001100011010111101110",
						 "100001100011011011101010",
						 "100001100011011111100110",
						 "100001100011100011100010",
						 "100001100011100111011110",
						 "100001100011101011011010",
						 "100001100011101111010110",
						 "100001100011110011010010",
						 "100001100011110111001110",
						 "100001100011111011001010",
						 "100001100011111111000110",
						 "100001100100000011000010",
						 "100001100100000110111110",
						 "100001100100001010111010",
						 "100001100100001110110110",
						 "100001100101110110110000",
						 "100001100101111010101100",
						 "100001100101111110101000",
						 "100001100110000010100100",
						 "100001100110000110100000",
						 "100001100110001010011100",
						 "100001100110001110011000",
						 "100001100110010010010100",
						 "100001100110010110010000",
						 "100001100110011010001100",
						 "100001100110011110001000",
						 "100001100110100010000100",
						 "100001100110100110000000",
						 "100001100110101001111100",
						 "100001100110101101111000",
						 "100001100110110001110100",
						 "100001100101110110110000",
						 "100001100101111010101100",
						 "100001100101111110101000",
						 "100001100110000010100100",
						 "100001100110000110100000",
						 "100001100110001010011100",
						 "100001100110001110011000",
						 "100001100110010010010100",
						 "100001100110010110010000",
						 "100001100110011010001100",
						 "100001100110011110001000",
						 "100001100110100010000100",
						 "100001100110100110000000",
						 "100001100110101001111100",
						 "100001100110101101111000",
						 "100001100110110001110100",
						 "100001101000011001101110",
						 "100001101000011101101010",
						 "100001101000100001100110",
						 "100001101000100101100010",
						 "100001101000101001011110",
						 "100001101000101101011010",
						 "100001101000110001010110",
						 "100001101000110101010010",
						 "100001101000111001001110",
						 "100001101000111101001010",
						 "100001101001000001000110",
						 "100001101001000101000010",
						 "100001101001001000111110",
						 "100001101001001100111010",
						 "100001101001010000110110",
						 "100001101001010100110010",
						 "100001101000011001101110",
						 "100001101000011101101010",
						 "100001101000100001100110",
						 "100001101000100101100010",
						 "100001101000101001011110",
						 "100001101000101101011010",
						 "100001101000110001010110",
						 "100001101000110101010010",
						 "100001101000111001001110",
						 "100001101000111101001010",
						 "100001101001000001000110",
						 "100001101001000101000010",
						 "100001101001001000111110",
						 "100001101001001100111010",
						 "100001101001010000110110",
						 "100001101001010100110010",
						 "100001101000011001101110",
						 "100001101000011101101010",
						 "100001101000100001100110",
						 "100001101000100101100010",
						 "100001101000101001011110",
						 "100001101000101101011010",
						 "100001101000110001010110",
						 "100001101000110101010010",
						 "100001101000111001001110",
						 "100001101000111101001010",
						 "100001101001000001000110",
						 "100001101001000101000010",
						 "100001101001001000111110",
						 "100001101001001100111010",
						 "100001101001010000110110",
						 "100001101001010100110010",
						 "100001101010111100101100",
						 "100001101011000000101000",
						 "100001101011000100100100",
						 "100001101011001000100000",
						 "100001101011001100011100",
						 "100001101011010000011000",
						 "100001101011010100010100",
						 "100001101011011000010000",
						 "100001101011011100001100",
						 "100001101011100000001000",
						 "100001101011100100000100",
						 "100001101011101000000000",
						 "100001101011101011111100",
						 "100001101011101111111000",
						 "100001101011110011110100",
						 "100001101011110111110000",
						 "100001101010111100101100",
						 "100001101011000000100111",
						 "100001101011000100100010",
						 "100001101011001000011101",
						 "100001101011001100011000",
						 "100001101011010000010011",
						 "100001101011010100001110",
						 "100001101011011000001001",
						 "100001101011011100000100",
						 "100001101011011111111111",
						 "100001101011100011111010",
						 "100001101011100111110101",
						 "100001101011101011110000",
						 "100001101011101111101011",
						 "100001101011110011100110",
						 "100001101011110111100001",
						 "100001101010111100101100",
						 "100001101011000000100111",
						 "100001101011000100100010",
						 "100001101011001000011101",
						 "100001101011001100011000",
						 "100001101011010000010011",
						 "100001101011010100001110",
						 "100001101011011000001001",
						 "100001101011011100000100",
						 "100001101011011111111111",
						 "100001101011100011111010",
						 "100001101011100111110101",
						 "100001101011101011110000",
						 "100001101011101111101011",
						 "100001101011110011100110",
						 "100001101011110111100001",
						 "100001101101011111101010",
						 "100001101101100011100101",
						 "100001101101100111100000",
						 "100001101101101011011011",
						 "100001101101101111010110",
						 "100001101101110011010001",
						 "100001101101110111001100",
						 "100001101101111011000111",
						 "100001101101111111000010",
						 "100001101110000010111101",
						 "100001101110000110111000",
						 "100001101110001010110011",
						 "100001101110001110101110",
						 "100001101110010010101001",
						 "100001101110010110100100",
						 "100001101110011010011111",
						 "100001101101011111101010",
						 "100001101101100011100101",
						 "100001101101100111100000",
						 "100001101101101011011011",
						 "100001101101101111010110",
						 "100001101101110011010001",
						 "100001101101110111001100",
						 "100001101101111011000111",
						 "100001101101111111000010",
						 "100001101110000010111101",
						 "100001101110000110111000",
						 "100001101110001010110011",
						 "100001101110001110101110",
						 "100001101110010010101001",
						 "100001101110010110100100",
						 "100001101110011010011111",
						 "100001110000000010101000",
						 "100001110000000110100011",
						 "100001110000001010011110",
						 "100001110000001110011001",
						 "100001110000010010010100",
						 "100001110000010110001111",
						 "100001110000011010001010",
						 "100001110000011110000101",
						 "100001110000100010000000",
						 "100001110000100101111011",
						 "100001110000101001110110",
						 "100001110000101101110001",
						 "100001110000110001101100",
						 "100001110000110101100111",
						 "100001110000111001100010",
						 "100001110000111101011101",
						 "100001110000000010101000",
						 "100001110000000110100011",
						 "100001110000001010011110",
						 "100001110000001110011001",
						 "100001110000010010010100",
						 "100001110000010110001111",
						 "100001110000011010001010",
						 "100001110000011110000101",
						 "100001110000100010000000",
						 "100001110000100101111011",
						 "100001110000101001110110",
						 "100001110000101101110001",
						 "100001110000110001101100",
						 "100001110000110101100111",
						 "100001110000111001100010",
						 "100001110000111101011101",
						 "100001110000000010101000",
						 "100001110000000110100011",
						 "100001110000001010011110",
						 "100001110000001110011001",
						 "100001110000010010010100",
						 "100001110000010110001111",
						 "100001110000011010001010",
						 "100001110000011110000101",
						 "100001110000100010000000",
						 "100001110000100101111011",
						 "100001110000101001110110",
						 "100001110000101101110001",
						 "100001110000110001101100",
						 "100001110000110101100111",
						 "100001110000111001100010",
						 "100001110000111101011101",
						 "100001110010100101100110",
						 "100001110010101001100001",
						 "100001110010101101011100",
						 "100001110010110001010111",
						 "100001110010110101010010",
						 "100001110010111001001101",
						 "100001110010111101001000",
						 "100001110011000001000011",
						 "100001110011000100111110",
						 "100001110011001000111001",
						 "100001110011001100110100",
						 "100001110011010000101111",
						 "100001110011010100101010",
						 "100001110011011000100101",
						 "100001110011011100100000",
						 "100001110011100000011011",
						 "100001110010100101100110",
						 "100001110010101001100001",
						 "100001110010101101011100",
						 "100001110010110001010111",
						 "100001110010110101010010",
						 "100001110010111001001101",
						 "100001110010111101001000",
						 "100001110011000001000011",
						 "100001110011000100111110",
						 "100001110011001000111001",
						 "100001110011001100110100",
						 "100001110011010000101111",
						 "100001110011010100101010",
						 "100001110011011000100101",
						 "100001110011011100100000",
						 "100001110011100000011011",
						 "100001110101001000100100",
						 "100001110101001100011111",
						 "100001110101010000011010",
						 "100001110101010100010101",
						 "100001110101011000010000",
						 "100001110101011100001011",
						 "100001110101100000000110",
						 "100001110101100100000001",
						 "100001110101100111111100",
						 "100001110101101011110111",
						 "100001110101101111110010",
						 "100001110101110011101101",
						 "100001110101110111101000",
						 "100001110101111011100011",
						 "100001110101111111011110",
						 "100001110110000011011001",
						 "100001110101001000100100",
						 "100001110101001100011111",
						 "100001110101010000011010",
						 "100001110101010100010101",
						 "100001110101011000010000",
						 "100001110101011100001011",
						 "100001110101100000000110",
						 "100001110101100100000001",
						 "100001110101100111111100",
						 "100001110101101011110111",
						 "100001110101101111110010",
						 "100001110101110011101101",
						 "100001110101110111101000",
						 "100001110101111011100011",
						 "100001110101111111011110",
						 "100001110110000011011001",
						 "100001110101001000100100",
						 "100001110101001100011111",
						 "100001110101010000011010",
						 "100001110101010100010101",
						 "100001110101011000010000",
						 "100001110101011100001011",
						 "100001110101100000000110",
						 "100001110101100100000001",
						 "100001110101100111111100",
						 "100001110101101011110111",
						 "100001110101101111110010",
						 "100001110101110011101101",
						 "100001110101110111101000",
						 "100001110101111011100011",
						 "100001110101111111011110",
						 "100001110110000011011001",
						 "100001110111101011100010",
						 "100001110111101111011101",
						 "100001110111110011011000",
						 "100001110111110111010011",
						 "100001110111111011001110",
						 "100001110111111111001001",
						 "100001111000000011000100",
						 "100001111000000110111111",
						 "100001111000001010111010",
						 "100001111000001110110101",
						 "100001111000010010110000",
						 "100001111000010110101011",
						 "100001111000011010100110",
						 "100001111000011110100001",
						 "100001111000100010011100",
						 "100001111000100110010111",
						 "100001110111101011100010",
						 "100001110111101111011101",
						 "100001110111110011011000",
						 "100001110111110111010011",
						 "100001110111111011001110",
						 "100001110111111111001001",
						 "100001111000000011000100",
						 "100001111000000110111111",
						 "100001111000001010111010",
						 "100001111000001110110101",
						 "100001111000010010110000",
						 "100001111000010110101011",
						 "100001111000011010100110",
						 "100001111000011110100001",
						 "100001111000100010011100",
						 "100001111000100110010111",
						 "100001110111101011100010",
						 "100001110111101111011101",
						 "100001110111110011011000",
						 "100001110111110111010011",
						 "100001110111111011001110",
						 "100001110111111111001001",
						 "100001111000000011000100",
						 "100001111000000110111111",
						 "100001111000001010111010",
						 "100001111000001110110101",
						 "100001111000010010110000",
						 "100001111000010110101011",
						 "100001111000011010100110",
						 "100001111000011110100001",
						 "100001111000100010011100",
						 "100001111000100110010111",
						 "100001111010001110100000",
						 "100001111010010010011010",
						 "100001111010010110010100",
						 "100001111010011010001110",
						 "100001111010011110001000",
						 "100001111010100010000010",
						 "100001111010100101111100",
						 "100001111010101001110110",
						 "100001111010101101110000",
						 "100001111010110001101010",
						 "100001111010110101100100",
						 "100001111010111001011110",
						 "100001111010111101011000",
						 "100001111011000001010010",
						 "100001111011000101001100",
						 "100001111011001001000110",
						 "100001111010001110100000",
						 "100001111010010010011010",
						 "100001111010010110010100",
						 "100001111010011010001110",
						 "100001111010011110001000",
						 "100001111010100010000010",
						 "100001111010100101111100",
						 "100001111010101001110110",
						 "100001111010101101110000",
						 "100001111010110001101010",
						 "100001111010110101100100",
						 "100001111010111001011110",
						 "100001111010111101011000",
						 "100001111011000001010010",
						 "100001111011000101001100",
						 "100001111011001001000110",
						 "100001111100110001011110",
						 "100001111100110101011000",
						 "100001111100111001010010",
						 "100001111100111101001100",
						 "100001111101000001000110",
						 "100001111101000101000000",
						 "100001111101001000111010",
						 "100001111101001100110100",
						 "100001111101010000101110",
						 "100001111101010100101000",
						 "100001111101011000100010",
						 "100001111101011100011100",
						 "100001111101100000010110",
						 "100001111101100100010000",
						 "100001111101101000001010",
						 "100001111101101100000100",
						 "100001111100110001011110",
						 "100001111100110101011000",
						 "100001111100111001010010",
						 "100001111100111101001100",
						 "100001111101000001000110",
						 "100001111101000101000000",
						 "100001111101001000111010",
						 "100001111101001100110100",
						 "100001111101010000101110",
						 "100001111101010100101000",
						 "100001111101011000100010",
						 "100001111101011100011100",
						 "100001111101100000010110",
						 "100001111101100100010000",
						 "100001111101101000001010",
						 "100001111101101100000100",
						 "100001111100110001011110",
						 "100001111100110101011000",
						 "100001111100111001010010",
						 "100001111100111101001100",
						 "100001111101000001000110",
						 "100001111101000101000000",
						 "100001111101001000111010",
						 "100001111101001100110100",
						 "100001111101010000101110",
						 "100001111101010100101000",
						 "100001111101011000100010",
						 "100001111101011100011100",
						 "100001111101100000010110",
						 "100001111101100100010000",
						 "100001111101101000001010",
						 "100001111101101100000100",
						 "100001111111010100011100",
						 "100001111111011000010110",
						 "100001111111011100010000",
						 "100001111111100000001010",
						 "100001111111100100000100",
						 "100001111111100111111110",
						 "100001111111101011111000",
						 "100001111111101111110010",
						 "100001111111110011101100",
						 "100001111111110111100110",
						 "100001111111111011100000",
						 "100001111111111111011010",
						 "100010000000000011010100",
						 "100010000000000111001110",
						 "100010000000001011001000",
						 "100010000000001111000010",
						 "100001111111010100011100",
						 "100001111111011000010110",
						 "100001111111011100010000",
						 "100001111111100000001010",
						 "100001111111100100000100",
						 "100001111111100111111110",
						 "100001111111101011111000",
						 "100001111111101111110010",
						 "100001111111110011101100",
						 "100001111111110111100110",
						 "100001111111111011100000",
						 "100001111111111111011010",
						 "100010000000000011010100",
						 "100010000000000111001110",
						 "100010000000001011001000",
						 "100010000000001111000010",
						 "100010000001110111011010",
						 "100010000001111011010100",
						 "100010000001111111001110",
						 "100010000010000011001000",
						 "100010000010000111000010",
						 "100010000010001010111100",
						 "100010000010001110110110",
						 "100010000010010010110000",
						 "100010000010010110101010",
						 "100010000010011010100100",
						 "100010000010011110011110",
						 "100010000010100010011000",
						 "100010000010100110010010",
						 "100010000010101010001100",
						 "100010000010101110000110",
						 "100010000010110010000000",
						 "100010000001110111011010",
						 "100010000001111011010100",
						 "100010000001111111001110",
						 "100010000010000011001000",
						 "100010000010000111000010",
						 "100010000010001010111100",
						 "100010000010001110110110",
						 "100010000010010010110000",
						 "100010000010010110101010",
						 "100010000010011010100100",
						 "100010000010011110011110",
						 "100010000010100010011000",
						 "100010000010100110010010",
						 "100010000010101010001100",
						 "100010000010101110000110",
						 "100010000010110010000000",
						 "100010000001110111011010",
						 "100010000001111011010100",
						 "100010000001111111001110",
						 "100010000010000011001000",
						 "100010000010000111000010",
						 "100010000010001010111100",
						 "100010000010001110110110",
						 "100010000010010010110000",
						 "100010000010010110101010",
						 "100010000010011010100100",
						 "100010000010011110011110",
						 "100010000010100010011000",
						 "100010000010100110010010",
						 "100010000010101010001100",
						 "100010000010101110000110",
						 "100010000010110010000000",
						 "100010000100011010011000",
						 "100010000100011110010010",
						 "100010000100100010001100",
						 "100010000100100110000110",
						 "100010000100101010000000",
						 "100010000100101101111010",
						 "100010000100110001110100",
						 "100010000100110101101110",
						 "100010000100111001101000",
						 "100010000100111101100010",
						 "100010000101000001011100",
						 "100010000101000101010110",
						 "100010000101001001010000",
						 "100010000101001101001010",
						 "100010000101010001000100",
						 "100010000101010100111110",
						 "100010000100011010011000",
						 "100010000100011110010010",
						 "100010000100100010001100",
						 "100010000100100110000110",
						 "100010000100101010000000",
						 "100010000100101101111010",
						 "100010000100110001110100",
						 "100010000100110101101110",
						 "100010000100111001101000",
						 "100010000100111101100010",
						 "100010000101000001011100",
						 "100010000101000101010110",
						 "100010000101001001010000",
						 "100010000101001101001010",
						 "100010000101010001000100",
						 "100010000101010100111110",
						 "100010000100011010011000",
						 "100010000100011110010010",
						 "100010000100100010001100",
						 "100010000100100110000110",
						 "100010000100101010000000",
						 "100010000100101101111010",
						 "100010000100110001110100",
						 "100010000100110101101110",
						 "100010000100111001101000",
						 "100010000100111101100010",
						 "100010000101000001011100",
						 "100010000101000101010110",
						 "100010000101001001010000",
						 "100010000101001101001010",
						 "100010000101010001000100",
						 "100010000101010100111110",
						 "100010000110111101010110",
						 "100010000111000001001111",
						 "100010000111000101001000",
						 "100010000111001001000001",
						 "100010000111001100111010",
						 "100010000111010000110011",
						 "100010000111010100101100",
						 "100010000111011000100101",
						 "100010000111011100011110",
						 "100010000111100000010111",
						 "100010000111100100010000",
						 "100010000111101000001001",
						 "100010000111101100000010",
						 "100010000111101111111011",
						 "100010000111110011110100",
						 "100010000111110111101101",
						 "100010000110111101010110",
						 "100010000111000001001111",
						 "100010000111000101001000",
						 "100010000111001001000001",
						 "100010000111001100111010",
						 "100010000111010000110011",
						 "100010000111010100101100",
						 "100010000111011000100101",
						 "100010000111011100011110",
						 "100010000111100000010111",
						 "100010000111100100010000",
						 "100010000111101000001001",
						 "100010000111101100000010",
						 "100010000111101111111011",
						 "100010000111110011110100",
						 "100010000111110111101101",
						 "100010001001100000010100",
						 "100010001001100100001101",
						 "100010001001101000000110",
						 "100010001001101011111111",
						 "100010001001101111111000",
						 "100010001001110011110001",
						 "100010001001110111101010",
						 "100010001001111011100011",
						 "100010001001111111011100",
						 "100010001010000011010101",
						 "100010001010000111001110",
						 "100010001010001011000111",
						 "100010001010001111000000",
						 "100010001010010010111001",
						 "100010001010010110110010",
						 "100010001010011010101011",
						 "100010001001100000010100",
						 "100010001001100100001101",
						 "100010001001101000000110",
						 "100010001001101011111111",
						 "100010001001101111111000",
						 "100010001001110011110001",
						 "100010001001110111101010",
						 "100010001001111011100011",
						 "100010001001111111011100",
						 "100010001010000011010101",
						 "100010001010000111001110",
						 "100010001010001011000111",
						 "100010001010001111000000",
						 "100010001010010010111001",
						 "100010001010010110110010",
						 "100010001010011010101011",
						 "100010001001100000010100",
						 "100010001001100100001101",
						 "100010001001101000000110",
						 "100010001001101011111111",
						 "100010001001101111111000",
						 "100010001001110011110001",
						 "100010001001110111101010",
						 "100010001001111011100011",
						 "100010001001111111011100",
						 "100010001010000011010101",
						 "100010001010000111001110",
						 "100010001010001011000111",
						 "100010001010001111000000",
						 "100010001010010010111001",
						 "100010001010010110110010",
						 "100010001010011010101011",
						 "100010001100000011010010",
						 "100010001100000111001011",
						 "100010001100001011000100",
						 "100010001100001110111101",
						 "100010001100010010110110",
						 "100010001100010110101111",
						 "100010001100011010101000",
						 "100010001100011110100001",
						 "100010001100100010011010",
						 "100010001100100110010011",
						 "100010001100101010001100",
						 "100010001100101110000101",
						 "100010001100110001111110",
						 "100010001100110101110111",
						 "100010001100111001110000",
						 "100010001100111101101001",
						 "100010001100000011010010",
						 "100010001100000111001011",
						 "100010001100001011000100",
						 "100010001100001110111101",
						 "100010001100010010110110",
						 "100010001100010110101111",
						 "100010001100011010101000",
						 "100010001100011110100001",
						 "100010001100100010011010",
						 "100010001100100110010011",
						 "100010001100101010001100",
						 "100010001100101110000101",
						 "100010001100110001111110",
						 "100010001100110101110111",
						 "100010001100111001110000",
						 "100010001100111101101001",
						 "100010001100000011010010",
						 "100010001100000111001011",
						 "100010001100001011000100",
						 "100010001100001110111101",
						 "100010001100010010110110",
						 "100010001100010110101111",
						 "100010001100011010101000",
						 "100010001100011110100001",
						 "100010001100100010011010",
						 "100010001100100110010011",
						 "100010001100101010001100",
						 "100010001100101110000101",
						 "100010001100110001111110",
						 "100010001100110101110111",
						 "100010001100111001110000",
						 "100010001100111101101001",
						 "100010001110100110010000",
						 "100010001110101010001001",
						 "100010001110101110000010",
						 "100010001110110001111011",
						 "100010001110110101110100",
						 "100010001110111001101101",
						 "100010001110111101100110",
						 "100010001111000001011111",
						 "100010001111000101011000",
						 "100010001111001001010001",
						 "100010001111001101001010",
						 "100010001111010001000011",
						 "100010001111010100111100",
						 "100010001111011000110101",
						 "100010001111011100101110",
						 "100010001111100000100111",
						 "100010001110100110010000",
						 "100010001110101010001001",
						 "100010001110101110000010",
						 "100010001110110001111011",
						 "100010001110110101110100",
						 "100010001110111001101101",
						 "100010001110111101100110",
						 "100010001111000001011111",
						 "100010001111000101011000",
						 "100010001111001001010001",
						 "100010001111001101001010",
						 "100010001111010001000011",
						 "100010001111010100111100",
						 "100010001111011000110101",
						 "100010001111011100101110",
						 "100010001111100000100111",
						 "100010010001001001001110",
						 "100010010001001101000111",
						 "100010010001010001000000",
						 "100010010001010100111001",
						 "100010010001011000110010",
						 "100010010001011100101011",
						 "100010010001100000100100",
						 "100010010001100100011101",
						 "100010010001101000010110",
						 "100010010001101100001111",
						 "100010010001110000001000",
						 "100010010001110100000001",
						 "100010010001110111111010",
						 "100010010001111011110011",
						 "100010010001111111101100",
						 "100010010010000011100101",
						 "100010010001001001001110",
						 "100010010001001101000111",
						 "100010010001010001000000",
						 "100010010001010100111001",
						 "100010010001011000110010",
						 "100010010001011100101011",
						 "100010010001100000100100",
						 "100010010001100100011101",
						 "100010010001101000010110",
						 "100010010001101100001111",
						 "100010010001110000001000",
						 "100010010001110100000001",
						 "100010010001110111111010",
						 "100010010001111011110011",
						 "100010010001111111101100",
						 "100010010010000011100101",
						 "100010010001001001001110",
						 "100010010001001101000110",
						 "100010010001010000111110",
						 "100010010001010100110110",
						 "100010010001011000101110",
						 "100010010001011100100110",
						 "100010010001100000011110",
						 "100010010001100100010110",
						 "100010010001101000001110",
						 "100010010001101100000110",
						 "100010010001101111111110",
						 "100010010001110011110110",
						 "100010010001110111101110",
						 "100010010001111011100110",
						 "100010010001111111011110",
						 "100010010010000011010110",
						 "100010010011101100001100",
						 "100010010011110000000100",
						 "100010010011110011111100",
						 "100010010011110111110100",
						 "100010010011111011101100",
						 "100010010011111111100100",
						 "100010010100000011011100",
						 "100010010100000111010100",
						 "100010010100001011001100",
						 "100010010100001111000100",
						 "100010010100010010111100",
						 "100010010100010110110100",
						 "100010010100011010101100",
						 "100010010100011110100100",
						 "100010010100100010011100",
						 "100010010100100110010100",
						 "100010010011101100001100",
						 "100010010011110000000100",
						 "100010010011110011111100",
						 "100010010011110111110100",
						 "100010010011111011101100",
						 "100010010011111111100100",
						 "100010010100000011011100",
						 "100010010100000111010100",
						 "100010010100001011001100",
						 "100010010100001111000100",
						 "100010010100010010111100",
						 "100010010100010110110100",
						 "100010010100011010101100",
						 "100010010100011110100100",
						 "100010010100100010011100",
						 "100010010100100110010100",
						 "100010010110001111001010",
						 "100010010110010011000010",
						 "100010010110010110111010",
						 "100010010110011010110010",
						 "100010010110011110101010",
						 "100010010110100010100010",
						 "100010010110100110011010",
						 "100010010110101010010010",
						 "100010010110101110001010",
						 "100010010110110010000010",
						 "100010010110110101111010",
						 "100010010110111001110010",
						 "100010010110111101101010",
						 "100010010111000001100010",
						 "100010010111000101011010",
						 "100010010111001001010010",
						 "100010010110001111001010",
						 "100010010110010011000010",
						 "100010010110010110111010",
						 "100010010110011010110010",
						 "100010010110011110101010",
						 "100010010110100010100010",
						 "100010010110100110011010",
						 "100010010110101010010010",
						 "100010010110101110001010",
						 "100010010110110010000010",
						 "100010010110110101111010",
						 "100010010110111001110010",
						 "100010010110111101101010",
						 "100010010111000001100010",
						 "100010010111000101011010",
						 "100010010111001001010010",
						 "100010010110001111001010",
						 "100010010110010011000010",
						 "100010010110010110111010",
						 "100010010110011010110010",
						 "100010010110011110101010",
						 "100010010110100010100010",
						 "100010010110100110011010",
						 "100010010110101010010010",
						 "100010010110101110001010",
						 "100010010110110010000010",
						 "100010010110110101111010",
						 "100010010110111001110010",
						 "100010010110111101101010",
						 "100010010111000001100010",
						 "100010010111000101011010",
						 "100010010111001001010010",
						 "100010011000110010001000",
						 "100010011000110110000000",
						 "100010011000111001111000",
						 "100010011000111101110000",
						 "100010011001000001101000",
						 "100010011001000101100000",
						 "100010011001001001011000",
						 "100010011001001101010000",
						 "100010011001010001001000",
						 "100010011001010101000000",
						 "100010011001011000111000",
						 "100010011001011100110000",
						 "100010011001100000101000",
						 "100010011001100100100000",
						 "100010011001101000011000",
						 "100010011001101100010000",
						 "100010011000110010001000",
						 "100010011000110110000000",
						 "100010011000111001111000",
						 "100010011000111101110000",
						 "100010011001000001101000",
						 "100010011001000101100000",
						 "100010011001001001011000",
						 "100010011001001101010000",
						 "100010011001010001001000",
						 "100010011001010101000000",
						 "100010011001011000111000",
						 "100010011001011100110000",
						 "100010011001100000101000",
						 "100010011001100100100000",
						 "100010011001101000011000",
						 "100010011001101100010000",
						 "100010011000110010001000",
						 "100010011000110110000000",
						 "100010011000111001111000",
						 "100010011000111101110000",
						 "100010011001000001101000",
						 "100010011001000101100000",
						 "100010011001001001011000",
						 "100010011001001101010000",
						 "100010011001010001001000",
						 "100010011001010101000000",
						 "100010011001011000111000",
						 "100010011001011100110000",
						 "100010011001100000101000",
						 "100010011001100100100000",
						 "100010011001101000011000",
						 "100010011001101100010000",
						 "100010011011010101000110",
						 "100010011011011000111110",
						 "100010011011011100110110",
						 "100010011011100000101110",
						 "100010011011100100100110",
						 "100010011011101000011110",
						 "100010011011101100010110",
						 "100010011011110000001110",
						 "100010011011110100000110",
						 "100010011011110111111110",
						 "100010011011111011110110",
						 "100010011011111111101110",
						 "100010011100000011100110",
						 "100010011100000111011110",
						 "100010011100001011010110",
						 "100010011100001111001110",
						 "100010011011010101000110",
						 "100010011011011000111101",
						 "100010011011011100110100",
						 "100010011011100000101011",
						 "100010011011100100100010",
						 "100010011011101000011001",
						 "100010011011101100010000",
						 "100010011011110000000111",
						 "100010011011110011111110",
						 "100010011011110111110101",
						 "100010011011111011101100",
						 "100010011011111111100011",
						 "100010011100000011011010",
						 "100010011100000111010001",
						 "100010011100001011001000",
						 "100010011100001110111111",
						 "100010011101111000000100",
						 "100010011101111011111011",
						 "100010011101111111110010",
						 "100010011110000011101001",
						 "100010011110000111100000",
						 "100010011110001011010111",
						 "100010011110001111001110",
						 "100010011110010011000101",
						 "100010011110010110111100",
						 "100010011110011010110011",
						 "100010011110011110101010",
						 "100010011110100010100001",
						 "100010011110100110011000",
						 "100010011110101010001111",
						 "100010011110101110000110",
						 "100010011110110001111101",
						 "100010011101111000000100",
						 "100010011101111011111011",
						 "100010011101111111110010",
						 "100010011110000011101001",
						 "100010011110000111100000",
						 "100010011110001011010111",
						 "100010011110001111001110",
						 "100010011110010011000101",
						 "100010011110010110111100",
						 "100010011110011010110011",
						 "100010011110011110101010",
						 "100010011110100010100001",
						 "100010011110100110011000",
						 "100010011110101010001111",
						 "100010011110101110000110",
						 "100010011110110001111101",
						 "100010011101111000000100",
						 "100010011101111011111011",
						 "100010011101111111110010",
						 "100010011110000011101001",
						 "100010011110000111100000",
						 "100010011110001011010111",
						 "100010011110001111001110",
						 "100010011110010011000101",
						 "100010011110010110111100",
						 "100010011110011010110011",
						 "100010011110011110101010",
						 "100010011110100010100001",
						 "100010011110100110011000",
						 "100010011110101010001111",
						 "100010011110101110000110",
						 "100010011110110001111101",
						 "100010100000011011000010",
						 "100010100000011110111001",
						 "100010100000100010110000",
						 "100010100000100110100111",
						 "100010100000101010011110",
						 "100010100000101110010101",
						 "100010100000110010001100",
						 "100010100000110110000011",
						 "100010100000111001111010",
						 "100010100000111101110001",
						 "100010100001000001101000",
						 "100010100001000101011111",
						 "100010100001001001010110",
						 "100010100001001101001101",
						 "100010100001010001000100",
						 "100010100001010100111011",
						 "100010100000011011000010",
						 "100010100000011110111001",
						 "100010100000100010110000",
						 "100010100000100110100111",
						 "100010100000101010011110",
						 "100010100000101110010101",
						 "100010100000110010001100",
						 "100010100000110110000011",
						 "100010100000111001111010",
						 "100010100000111101110001",
						 "100010100001000001101000",
						 "100010100001000101011111",
						 "100010100001001001010110",
						 "100010100001001101001101",
						 "100010100001010001000100",
						 "100010100001010100111011",
						 "100010100000011011000010",
						 "100010100000011110111001",
						 "100010100000100010110000",
						 "100010100000100110100111",
						 "100010100000101010011110",
						 "100010100000101110010101",
						 "100010100000110010001100",
						 "100010100000110110000011",
						 "100010100000111001111010",
						 "100010100000111101110001",
						 "100010100001000001101000",
						 "100010100001000101011111",
						 "100010100001001001010110",
						 "100010100001001101001101",
						 "100010100001010001000100",
						 "100010100001010100111011",
						 "100010100010111110000000",
						 "100010100011000001110111",
						 "100010100011000101101110",
						 "100010100011001001100101",
						 "100010100011001101011100",
						 "100010100011010001010011",
						 "100010100011010101001010",
						 "100010100011011001000001",
						 "100010100011011100111000",
						 "100010100011100000101111",
						 "100010100011100100100110",
						 "100010100011101000011101",
						 "100010100011101100010100",
						 "100010100011110000001011",
						 "100010100011110100000010",
						 "100010100011110111111001",
						 "100010100010111110000000",
						 "100010100011000001110111",
						 "100010100011000101101110",
						 "100010100011001001100101",
						 "100010100011001101011100",
						 "100010100011010001010011",
						 "100010100011010101001010",
						 "100010100011011001000001",
						 "100010100011011100111000",
						 "100010100011100000101111",
						 "100010100011100100100110",
						 "100010100011101000011101",
						 "100010100011101100010100",
						 "100010100011110000001011",
						 "100010100011110100000010",
						 "100010100011110111111001",
						 "100010100101100000111110",
						 "100010100101100100110101",
						 "100010100101101000101100",
						 "100010100101101100100011",
						 "100010100101110000011010",
						 "100010100101110100010001",
						 "100010100101111000001000",
						 "100010100101111011111111",
						 "100010100101111111110110",
						 "100010100110000011101101",
						 "100010100110000111100100",
						 "100010100110001011011011",
						 "100010100110001111010010",
						 "100010100110010011001001",
						 "100010100110010111000000",
						 "100010100110011010110111",
						 "100010100101100000111110",
						 "100010100101100100110101",
						 "100010100101101000101100",
						 "100010100101101100100011",
						 "100010100101110000011010",
						 "100010100101110100010001",
						 "100010100101111000001000",
						 "100010100101111011111111",
						 "100010100101111111110110",
						 "100010100110000011101101",
						 "100010100110000111100100",
						 "100010100110001011011011",
						 "100010100110001111010010",
						 "100010100110010011001001",
						 "100010100110010111000000",
						 "100010100110011010110111",
						 "100010100101100000111110",
						 "100010100101100100110100",
						 "100010100101101000101010",
						 "100010100101101100100000",
						 "100010100101110000010110",
						 "100010100101110100001100",
						 "100010100101111000000010",
						 "100010100101111011111000",
						 "100010100101111111101110",
						 "100010100110000011100100",
						 "100010100110000111011010",
						 "100010100110001011010000",
						 "100010100110001111000110",
						 "100010100110010010111100",
						 "100010100110010110110010",
						 "100010100110011010101000",
						 "100010101000000011111100",
						 "100010101000000111110010",
						 "100010101000001011101000",
						 "100010101000001111011110",
						 "100010101000010011010100",
						 "100010101000010111001010",
						 "100010101000011011000000",
						 "100010101000011110110110",
						 "100010101000100010101100",
						 "100010101000100110100010",
						 "100010101000101010011000",
						 "100010101000101110001110",
						 "100010101000110010000100",
						 "100010101000110101111010",
						 "100010101000111001110000",
						 "100010101000111101100110",
						 "100010101000000011111100",
						 "100010101000000111110010",
						 "100010101000001011101000",
						 "100010101000001111011110",
						 "100010101000010011010100",
						 "100010101000010111001010",
						 "100010101000011011000000",
						 "100010101000011110110110",
						 "100010101000100010101100",
						 "100010101000100110100010",
						 "100010101000101010011000",
						 "100010101000101110001110",
						 "100010101000110010000100",
						 "100010101000110101111010",
						 "100010101000111001110000",
						 "100010101000111101100110",
						 "100010101010100110111010",
						 "100010101010101010110000",
						 "100010101010101110100110",
						 "100010101010110010011100",
						 "100010101010110110010010",
						 "100010101010111010001000",
						 "100010101010111101111110",
						 "100010101011000001110100",
						 "100010101011000101101010",
						 "100010101011001001100000",
						 "100010101011001101010110",
						 "100010101011010001001100",
						 "100010101011010101000010",
						 "100010101011011000111000",
						 "100010101011011100101110",
						 "100010101011100000100100",
						 "100010101010100110111010",
						 "100010101010101010110000",
						 "100010101010101110100110",
						 "100010101010110010011100",
						 "100010101010110110010010",
						 "100010101010111010001000",
						 "100010101010111101111110",
						 "100010101011000001110100",
						 "100010101011000101101010",
						 "100010101011001001100000",
						 "100010101011001101010110",
						 "100010101011010001001100",
						 "100010101011010101000010",
						 "100010101011011000111000",
						 "100010101011011100101110",
						 "100010101011100000100100",
						 "100010101010100110111010",
						 "100010101010101010110000",
						 "100010101010101110100110",
						 "100010101010110010011100",
						 "100010101010110110010010",
						 "100010101010111010001000",
						 "100010101010111101111110",
						 "100010101011000001110100",
						 "100010101011000101101010",
						 "100010101011001001100000",
						 "100010101011001101010110",
						 "100010101011010001001100",
						 "100010101011010101000010",
						 "100010101011011000111000",
						 "100010101011011100101110",
						 "100010101011100000100100",
						 "100010101101001001111000",
						 "100010101101001101101110",
						 "100010101101010001100100",
						 "100010101101010101011010",
						 "100010101101011001010000",
						 "100010101101011101000110",
						 "100010101101100000111100",
						 "100010101101100100110010",
						 "100010101101101000101000",
						 "100010101101101100011110",
						 "100010101101110000010100",
						 "100010101101110100001010",
						 "100010101101111000000000",
						 "100010101101111011110110",
						 "100010101101111111101100",
						 "100010101110000011100010",
						 "100010101101001001111000",
						 "100010101101001101101110",
						 "100010101101010001100100",
						 "100010101101010101011010",
						 "100010101101011001010000",
						 "100010101101011101000110",
						 "100010101101100000111100",
						 "100010101101100100110010",
						 "100010101101101000101000",
						 "100010101101101100011110",
						 "100010101101110000010100",
						 "100010101101110100001010",
						 "100010101101111000000000",
						 "100010101101111011110110",
						 "100010101101111111101100",
						 "100010101110000011100010",
						 "100010101101001001111000",
						 "100010101101001101101110",
						 "100010101101010001100100",
						 "100010101101010101011010",
						 "100010101101011001010000",
						 "100010101101011101000110",
						 "100010101101100000111100",
						 "100010101101100100110010",
						 "100010101101101000101000",
						 "100010101101101100011110",
						 "100010101101110000010100",
						 "100010101101110100001010",
						 "100010101101111000000000",
						 "100010101101111011110110",
						 "100010101101111111101100",
						 "100010101110000011100010",
						 "100010101111101100110110",
						 "100010101111110000101011",
						 "100010101111110100100000",
						 "100010101111111000010101",
						 "100010101111111100001010",
						 "100010101111111111111111",
						 "100010110000000011110100",
						 "100010110000000111101001",
						 "100010110000001011011110",
						 "100010110000001111010011",
						 "100010110000010011001000",
						 "100010110000010110111101",
						 "100010110000011010110010",
						 "100010110000011110100111",
						 "100010110000100010011100",
						 "100010110000100110010001",
						 "100010101111101100110110",
						 "100010101111110000101011",
						 "100010101111110100100000",
						 "100010101111111000010101",
						 "100010101111111100001010",
						 "100010101111111111111111",
						 "100010110000000011110100",
						 "100010110000000111101001",
						 "100010110000001011011110",
						 "100010110000001111010011",
						 "100010110000010011001000",
						 "100010110000010110111101",
						 "100010110000011010110010",
						 "100010110000011110100111",
						 "100010110000100010011100",
						 "100010110000100110010001",
						 "100010110010001111110100",
						 "100010110010010011101001",
						 "100010110010010111011110",
						 "100010110010011011010011",
						 "100010110010011111001000",
						 "100010110010100010111101",
						 "100010110010100110110010",
						 "100010110010101010100111",
						 "100010110010101110011100",
						 "100010110010110010010001",
						 "100010110010110110000110",
						 "100010110010111001111011",
						 "100010110010111101110000",
						 "100010110011000001100101",
						 "100010110011000101011010",
						 "100010110011001001001111",
						 "100010110010001111110100",
						 "100010110010010011101001",
						 "100010110010010111011110",
						 "100010110010011011010011",
						 "100010110010011111001000",
						 "100010110010100010111101",
						 "100010110010100110110010",
						 "100010110010101010100111",
						 "100010110010101110011100",
						 "100010110010110010010001",
						 "100010110010110110000110",
						 "100010110010111001111011",
						 "100010110010111101110000",
						 "100010110011000001100101",
						 "100010110011000101011010",
						 "100010110011001001001111",
						 "100010110010001111110100",
						 "100010110010010011101001",
						 "100010110010010111011110",
						 "100010110010011011010011",
						 "100010110010011111001000",
						 "100010110010100010111101",
						 "100010110010100110110010",
						 "100010110010101010100111",
						 "100010110010101110011100",
						 "100010110010110010010001",
						 "100010110010110110000110",
						 "100010110010111001111011",
						 "100010110010111101110000",
						 "100010110011000001100101",
						 "100010110011000101011010",
						 "100010110011001001001111",
						 "100010110100110010110010",
						 "100010110100110110100111",
						 "100010110100111010011100",
						 "100010110100111110010001",
						 "100010110101000010000110",
						 "100010110101000101111011",
						 "100010110101001001110000",
						 "100010110101001101100101",
						 "100010110101010001011010",
						 "100010110101010101001111",
						 "100010110101011001000100",
						 "100010110101011100111001",
						 "100010110101100000101110",
						 "100010110101100100100011",
						 "100010110101101000011000",
						 "100010110101101100001101",
						 "100010110100110010110010",
						 "100010110100110110100111",
						 "100010110100111010011100",
						 "100010110100111110010001",
						 "100010110101000010000110",
						 "100010110101000101111011",
						 "100010110101001001110000",
						 "100010110101001101100101",
						 "100010110101010001011010",
						 "100010110101010101001111",
						 "100010110101011001000100",
						 "100010110101011100111001",
						 "100010110101100000101110",
						 "100010110101100100100011",
						 "100010110101101000011000",
						 "100010110101101100001101",
						 "100010110100110010110010",
						 "100010110100110110100111",
						 "100010110100111010011100",
						 "100010110100111110010001",
						 "100010110101000010000110",
						 "100010110101000101111011",
						 "100010110101001001110000",
						 "100010110101001101100101",
						 "100010110101010001011010",
						 "100010110101010101001111",
						 "100010110101011001000100",
						 "100010110101011100111001",
						 "100010110101100000101110",
						 "100010110101100100100011",
						 "100010110101101000011000",
						 "100010110101101100001101",
						 "100010110111010101110000",
						 "100010110111011001100101",
						 "100010110111011101011010",
						 "100010110111100001001111",
						 "100010110111100101000100",
						 "100010110111101000111001",
						 "100010110111101100101110",
						 "100010110111110000100011",
						 "100010110111110100011000",
						 "100010110111111000001101",
						 "100010110111111100000010",
						 "100010110111111111110111",
						 "100010111000000011101100",
						 "100010111000000111100001",
						 "100010111000001011010110",
						 "100010111000001111001011",
						 "100010110111010101110000",
						 "100010110111011001100101",
						 "100010110111011101011010",
						 "100010110111100001001111",
						 "100010110111100101000100",
						 "100010110111101000111001",
						 "100010110111101100101110",
						 "100010110111110000100011",
						 "100010110111110100011000",
						 "100010110111111000001101",
						 "100010110111111100000010",
						 "100010110111111111110111",
						 "100010111000000011101100",
						 "100010111000000111100001",
						 "100010111000001011010110",
						 "100010111000001111001011",
						 "100010111001111000101110",
						 "100010111001111100100010",
						 "100010111010000000010110",
						 "100010111010000100001010",
						 "100010111010000111111110",
						 "100010111010001011110010",
						 "100010111010001111100110",
						 "100010111010010011011010",
						 "100010111010010111001110",
						 "100010111010011011000010",
						 "100010111010011110110110",
						 "100010111010100010101010",
						 "100010111010100110011110",
						 "100010111010101010010010",
						 "100010111010101110000110",
						 "100010111010110001111010",
						 "100010111001111000101110",
						 "100010111001111100100010",
						 "100010111010000000010110",
						 "100010111010000100001010",
						 "100010111010000111111110",
						 "100010111010001011110010",
						 "100010111010001111100110",
						 "100010111010010011011010",
						 "100010111010010111001110",
						 "100010111010011011000010",
						 "100010111010011110110110",
						 "100010111010100010101010",
						 "100010111010100110011110",
						 "100010111010101010010010",
						 "100010111010101110000110",
						 "100010111010110001111010",
						 "100010111001111000101110",
						 "100010111001111100100010",
						 "100010111010000000010110",
						 "100010111010000100001010",
						 "100010111010000111111110",
						 "100010111010001011110010",
						 "100010111010001111100110",
						 "100010111010010011011010",
						 "100010111010010111001110",
						 "100010111010011011000010",
						 "100010111010011110110110",
						 "100010111010100010101010",
						 "100010111010100110011110",
						 "100010111010101010010010",
						 "100010111010101110000110",
						 "100010111010110001111010",
						 "100010111100011011101100",
						 "100010111100011111100000",
						 "100010111100100011010100",
						 "100010111100100111001000",
						 "100010111100101010111100",
						 "100010111100101110110000",
						 "100010111100110010100100",
						 "100010111100110110011000",
						 "100010111100111010001100",
						 "100010111100111110000000",
						 "100010111101000001110100",
						 "100010111101000101101000",
						 "100010111101001001011100",
						 "100010111101001101010000",
						 "100010111101010001000100",
						 "100010111101010100111000",
						 "100010111100011011101100",
						 "100010111100011111100000",
						 "100010111100100011010100",
						 "100010111100100111001000",
						 "100010111100101010111100",
						 "100010111100101110110000",
						 "100010111100110010100100",
						 "100010111100110110011000",
						 "100010111100111010001100",
						 "100010111100111110000000",
						 "100010111101000001110100",
						 "100010111101000101101000",
						 "100010111101001001011100",
						 "100010111101001101010000",
						 "100010111101010001000100",
						 "100010111101010100111000",
						 "100010111100011011101100",
						 "100010111100011111100000",
						 "100010111100100011010100",
						 "100010111100100111001000",
						 "100010111100101010111100",
						 "100010111100101110110000",
						 "100010111100110010100100",
						 "100010111100110110011000",
						 "100010111100111010001100",
						 "100010111100111110000000",
						 "100010111101000001110100",
						 "100010111101000101101000",
						 "100010111101001001011100",
						 "100010111101001101010000",
						 "100010111101010001000100",
						 "100010111101010100111000",
						 "100010111110111110101010",
						 "100010111111000010011110",
						 "100010111111000110010010",
						 "100010111111001010000110",
						 "100010111111001101111010",
						 "100010111111010001101110",
						 "100010111111010101100010",
						 "100010111111011001010110",
						 "100010111111011101001010",
						 "100010111111100000111110",
						 "100010111111100100110010",
						 "100010111111101000100110",
						 "100010111111101100011010",
						 "100010111111110000001110",
						 "100010111111110100000010",
						 "100010111111110111110110",
						 "100010111110111110101010",
						 "100010111111000010011110",
						 "100010111111000110010010",
						 "100010111111001010000110",
						 "100010111111001101111010",
						 "100010111111010001101110",
						 "100010111111010101100010",
						 "100010111111011001010110",
						 "100010111111011101001010",
						 "100010111111100000111110",
						 "100010111111100100110010",
						 "100010111111101000100110",
						 "100010111111101100011010",
						 "100010111111110000001110",
						 "100010111111110100000010",
						 "100010111111110111110110",
						 "100011000001100001101000",
						 "100011000001100101011100",
						 "100011000001101001010000",
						 "100011000001101101000100",
						 "100011000001110000111000",
						 "100011000001110100101100",
						 "100011000001111000100000",
						 "100011000001111100010100",
						 "100011000010000000001000",
						 "100011000010000011111100",
						 "100011000010000111110000",
						 "100011000010001011100100",
						 "100011000010001111011000",
						 "100011000010010011001100",
						 "100011000010010111000000",
						 "100011000010011010110100",
						 "100011000001100001101000",
						 "100011000001100101011011",
						 "100011000001101001001110",
						 "100011000001101101000001",
						 "100011000001110000110100",
						 "100011000001110100100111",
						 "100011000001111000011010",
						 "100011000001111100001101",
						 "100011000010000000000000",
						 "100011000010000011110011",
						 "100011000010000111100110",
						 "100011000010001011011001",
						 "100011000010001111001100",
						 "100011000010010010111111",
						 "100011000010010110110010",
						 "100011000010011010100101",
						 "100011000001100001101000",
						 "100011000001100101011011",
						 "100011000001101001001110",
						 "100011000001101101000001",
						 "100011000001110000110100",
						 "100011000001110100100111",
						 "100011000001111000011010",
						 "100011000001111100001101",
						 "100011000010000000000000",
						 "100011000010000011110011",
						 "100011000010000111100110",
						 "100011000010001011011001",
						 "100011000010001111001100",
						 "100011000010010010111111",
						 "100011000010010110110010",
						 "100011000010011010100101",
						 "100011000100000100100110",
						 "100011000100001000011001",
						 "100011000100001100001100",
						 "100011000100001111111111",
						 "100011000100010011110010",
						 "100011000100010111100101",
						 "100011000100011011011000",
						 "100011000100011111001011",
						 "100011000100100010111110",
						 "100011000100100110110001",
						 "100011000100101010100100",
						 "100011000100101110010111",
						 "100011000100110010001010",
						 "100011000100110101111101",
						 "100011000100111001110000",
						 "100011000100111101100011",
						 "100011000100000100100110",
						 "100011000100001000011001",
						 "100011000100001100001100",
						 "100011000100001111111111",
						 "100011000100010011110010",
						 "100011000100010111100101",
						 "100011000100011011011000",
						 "100011000100011111001011",
						 "100011000100100010111110",
						 "100011000100100110110001",
						 "100011000100101010100100",
						 "100011000100101110010111",
						 "100011000100110010001010",
						 "100011000100110101111101",
						 "100011000100111001110000",
						 "100011000100111101100011",
						 "100011000100000100100110",
						 "100011000100001000011001",
						 "100011000100001100001100",
						 "100011000100001111111111",
						 "100011000100010011110010",
						 "100011000100010111100101",
						 "100011000100011011011000",
						 "100011000100011111001011",
						 "100011000100100010111110",
						 "100011000100100110110001",
						 "100011000100101010100100",
						 "100011000100101110010111",
						 "100011000100110010001010",
						 "100011000100110101111101",
						 "100011000100111001110000",
						 "100011000100111101100011",
						 "100011000110100111100100",
						 "100011000110101011010111",
						 "100011000110101111001010",
						 "100011000110110010111101",
						 "100011000110110110110000",
						 "100011000110111010100011",
						 "100011000110111110010110",
						 "100011000111000010001001",
						 "100011000111000101111100",
						 "100011000111001001101111",
						 "100011000111001101100010",
						 "100011000111010001010101",
						 "100011000111010101001000",
						 "100011000111011000111011",
						 "100011000111011100101110",
						 "100011000111100000100001",
						 "100011000110100111100100",
						 "100011000110101011010111",
						 "100011000110101111001010",
						 "100011000110110010111101",
						 "100011000110110110110000",
						 "100011000110111010100011",
						 "100011000110111110010110",
						 "100011000111000010001001",
						 "100011000111000101111100",
						 "100011000111001001101111",
						 "100011000111001101100010",
						 "100011000111010001010101",
						 "100011000111010101001000",
						 "100011000111011000111011",
						 "100011000111011100101110",
						 "100011000111100000100001",
						 "100011001001001010100010",
						 "100011001001001110010101",
						 "100011001001010010001000",
						 "100011001001010101111011",
						 "100011001001011001101110",
						 "100011001001011101100001",
						 "100011001001100001010100",
						 "100011001001100101000111",
						 "100011001001101000111010",
						 "100011001001101100101101",
						 "100011001001110000100000",
						 "100011001001110100010011",
						 "100011001001111000000110",
						 "100011001001111011111001",
						 "100011001001111111101100",
						 "100011001010000011011111",
						 "100011001001001010100010",
						 "100011001001001110010100",
						 "100011001001010010000110",
						 "100011001001010101111000",
						 "100011001001011001101010",
						 "100011001001011101011100",
						 "100011001001100001001110",
						 "100011001001100101000000",
						 "100011001001101000110010",
						 "100011001001101100100100",
						 "100011001001110000010110",
						 "100011001001110100001000",
						 "100011001001110111111010",
						 "100011001001111011101100",
						 "100011001001111111011110",
						 "100011001010000011010000",
						 "100011001001001010100010",
						 "100011001001001110010100",
						 "100011001001010010000110",
						 "100011001001010101111000",
						 "100011001001011001101010",
						 "100011001001011101011100",
						 "100011001001100001001110",
						 "100011001001100101000000",
						 "100011001001101000110010",
						 "100011001001101100100100",
						 "100011001001110000010110",
						 "100011001001110100001000",
						 "100011001001110111111010",
						 "100011001001111011101100",
						 "100011001001111111011110",
						 "100011001010000011010000",
						 "100011001011101101100000",
						 "100011001011110001010010",
						 "100011001011110101000100",
						 "100011001011111000110110",
						 "100011001011111100101000",
						 "100011001100000000011010",
						 "100011001100000100001100",
						 "100011001100000111111110",
						 "100011001100001011110000",
						 "100011001100001111100010",
						 "100011001100010011010100",
						 "100011001100010111000110",
						 "100011001100011010111000",
						 "100011001100011110101010",
						 "100011001100100010011100",
						 "100011001100100110001110",
						 "100011001011101101100000",
						 "100011001011110001010010",
						 "100011001011110101000100",
						 "100011001011111000110110",
						 "100011001011111100101000",
						 "100011001100000000011010",
						 "100011001100000100001100",
						 "100011001100000111111110",
						 "100011001100001011110000",
						 "100011001100001111100010",
						 "100011001100010011010100",
						 "100011001100010111000110",
						 "100011001100011010111000",
						 "100011001100011110101010",
						 "100011001100100010011100",
						 "100011001100100110001110",
						 "100011001011101101100000",
						 "100011001011110001010010",
						 "100011001011110101000100",
						 "100011001011111000110110",
						 "100011001011111100101000",
						 "100011001100000000011010",
						 "100011001100000100001100",
						 "100011001100000111111110",
						 "100011001100001011110000",
						 "100011001100001111100010",
						 "100011001100010011010100",
						 "100011001100010111000110",
						 "100011001100011010111000",
						 "100011001100011110101010",
						 "100011001100100010011100",
						 "100011001100100110001110",
						 "100011001110010000011110",
						 "100011001110010100010000",
						 "100011001110011000000010",
						 "100011001110011011110100",
						 "100011001110011111100110",
						 "100011001110100011011000",
						 "100011001110100111001010",
						 "100011001110101010111100",
						 "100011001110101110101110",
						 "100011001110110010100000",
						 "100011001110110110010010",
						 "100011001110111010000100",
						 "100011001110111101110110",
						 "100011001111000001101000",
						 "100011001111000101011010",
						 "100011001111001001001100",
						 "100011001110010000011110",
						 "100011001110010100010000",
						 "100011001110011000000010",
						 "100011001110011011110100",
						 "100011001110011111100110",
						 "100011001110100011011000",
						 "100011001110100111001010",
						 "100011001110101010111100",
						 "100011001110101110101110",
						 "100011001110110010100000",
						 "100011001110110110010010",
						 "100011001110111010000100",
						 "100011001110111101110110",
						 "100011001111000001101000",
						 "100011001111000101011010",
						 "100011001111001001001100",
						 "100011001110010000011110",
						 "100011001110010100010000",
						 "100011001110011000000010",
						 "100011001110011011110100",
						 "100011001110011111100110",
						 "100011001110100011011000",
						 "100011001110100111001010",
						 "100011001110101010111100",
						 "100011001110101110101110",
						 "100011001110110010100000",
						 "100011001110110110010010",
						 "100011001110111010000100",
						 "100011001110111101110110",
						 "100011001111000001101000",
						 "100011001111000101011010",
						 "100011001111001001001100",
						 "100011010000110011011100",
						 "100011010000110111001101",
						 "100011010000111010111110",
						 "100011010000111110101111",
						 "100011010001000010100000",
						 "100011010001000110010001",
						 "100011010001001010000010",
						 "100011010001001101110011",
						 "100011010001010001100100",
						 "100011010001010101010101",
						 "100011010001011001000110",
						 "100011010001011100110111",
						 "100011010001100000101000",
						 "100011010001100100011001",
						 "100011010001101000001010",
						 "100011010001101011111011",
						 "100011010000110011011100",
						 "100011010000110111001101",
						 "100011010000111010111110",
						 "100011010000111110101111",
						 "100011010001000010100000",
						 "100011010001000110010001",
						 "100011010001001010000010",
						 "100011010001001101110011",
						 "100011010001010001100100",
						 "100011010001010101010101",
						 "100011010001011001000110",
						 "100011010001011100110111",
						 "100011010001100000101000",
						 "100011010001100100011001",
						 "100011010001101000001010",
						 "100011010001101011111011",
						 "100011010011010110011010",
						 "100011010011011010001011",
						 "100011010011011101111100",
						 "100011010011100001101101",
						 "100011010011100101011110",
						 "100011010011101001001111",
						 "100011010011101101000000",
						 "100011010011110000110001",
						 "100011010011110100100010",
						 "100011010011111000010011",
						 "100011010011111100000100",
						 "100011010011111111110101",
						 "100011010100000011100110",
						 "100011010100000111010111",
						 "100011010100001011001000",
						 "100011010100001110111001",
						 "100011010011010110011010",
						 "100011010011011010001011",
						 "100011010011011101111100",
						 "100011010011100001101101",
						 "100011010011100101011110",
						 "100011010011101001001111",
						 "100011010011101101000000",
						 "100011010011110000110001",
						 "100011010011110100100010",
						 "100011010011111000010011",
						 "100011010011111100000100",
						 "100011010011111111110101",
						 "100011010100000011100110",
						 "100011010100000111010111",
						 "100011010100001011001000",
						 "100011010100001110111001",
						 "100011010011010110011010",
						 "100011010011011010001011",
						 "100011010011011101111100",
						 "100011010011100001101101",
						 "100011010011100101011110",
						 "100011010011101001001111",
						 "100011010011101101000000",
						 "100011010011110000110001",
						 "100011010011110100100010",
						 "100011010011111000010011",
						 "100011010011111100000100",
						 "100011010011111111110101",
						 "100011010100000011100110",
						 "100011010100000111010111",
						 "100011010100001011001000",
						 "100011010100001110111001",
						 "100011010101111001011000",
						 "100011010101111101001001",
						 "100011010110000000111010",
						 "100011010110000100101011",
						 "100011010110001000011100",
						 "100011010110001100001101",
						 "100011010110001111111110",
						 "100011010110010011101111",
						 "100011010110010111100000",
						 "100011010110011011010001",
						 "100011010110011111000010",
						 "100011010110100010110011",
						 "100011010110100110100100",
						 "100011010110101010010101",
						 "100011010110101110000110",
						 "100011010110110001110111",
						 "100011010101111001011000",
						 "100011010101111101001001",
						 "100011010110000000111010",
						 "100011010110000100101011",
						 "100011010110001000011100",
						 "100011010110001100001101",
						 "100011010110001111111110",
						 "100011010110010011101111",
						 "100011010110010111100000",
						 "100011010110011011010001",
						 "100011010110011111000010",
						 "100011010110100010110011",
						 "100011010110100110100100",
						 "100011010110101010010101",
						 "100011010110101110000110",
						 "100011010110110001110111",
						 "100011010101111001011000",
						 "100011010101111101001001",
						 "100011010110000000111010",
						 "100011010110000100101011",
						 "100011010110001000011100",
						 "100011010110001100001101",
						 "100011010110001111111110",
						 "100011010110010011101111",
						 "100011010110010111100000",
						 "100011010110011011010001",
						 "100011010110011111000010",
						 "100011010110100010110011",
						 "100011010110100110100100",
						 "100011010110101010010101",
						 "100011010110101110000110",
						 "100011010110110001110111",
						 "100011011000011100010110",
						 "100011011000100000000110",
						 "100011011000100011110110",
						 "100011011000100111100110",
						 "100011011000101011010110",
						 "100011011000101111000110",
						 "100011011000110010110110",
						 "100011011000110110100110",
						 "100011011000111010010110",
						 "100011011000111110000110",
						 "100011011001000001110110",
						 "100011011001000101100110",
						 "100011011001001001010110",
						 "100011011001001101000110",
						 "100011011001010000110110",
						 "100011011001010100100110",
						 "100011011000011100010110",
						 "100011011000100000000110",
						 "100011011000100011110110",
						 "100011011000100111100110",
						 "100011011000101011010110",
						 "100011011000101111000110",
						 "100011011000110010110110",
						 "100011011000110110100110",
						 "100011011000111010010110",
						 "100011011000111110000110",
						 "100011011001000001110110",
						 "100011011001000101100110",
						 "100011011001001001010110",
						 "100011011001001101000110",
						 "100011011001010000110110",
						 "100011011001010100100110",
						 "100011011010111111010100",
						 "100011011011000011000100",
						 "100011011011000110110100",
						 "100011011011001010100100",
						 "100011011011001110010100",
						 "100011011011010010000100",
						 "100011011011010101110100",
						 "100011011011011001100100",
						 "100011011011011101010100",
						 "100011011011100001000100",
						 "100011011011100100110100",
						 "100011011011101000100100",
						 "100011011011101100010100",
						 "100011011011110000000100",
						 "100011011011110011110100",
						 "100011011011110111100100",
						 "100011011010111111010100",
						 "100011011011000011000100",
						 "100011011011000110110100",
						 "100011011011001010100100",
						 "100011011011001110010100",
						 "100011011011010010000100",
						 "100011011011010101110100",
						 "100011011011011001100100",
						 "100011011011011101010100",
						 "100011011011100001000100",
						 "100011011011100100110100",
						 "100011011011101000100100",
						 "100011011011101100010100",
						 "100011011011110000000100",
						 "100011011011110011110100",
						 "100011011011110111100100",
						 "100011011010111111010100",
						 "100011011011000011000100",
						 "100011011011000110110100",
						 "100011011011001010100100",
						 "100011011011001110010100",
						 "100011011011010010000100",
						 "100011011011010101110100",
						 "100011011011011001100100",
						 "100011011011011101010100",
						 "100011011011100001000100",
						 "100011011011100100110100",
						 "100011011011101000100100",
						 "100011011011101100010100",
						 "100011011011110000000100",
						 "100011011011110011110100",
						 "100011011011110111100100",
						 "100011011101100010010010",
						 "100011011101100110000010",
						 "100011011101101001110010",
						 "100011011101101101100010",
						 "100011011101110001010010",
						 "100011011101110101000010",
						 "100011011101111000110010",
						 "100011011101111100100010",
						 "100011011110000000010010",
						 "100011011110000100000010",
						 "100011011110000111110010",
						 "100011011110001011100010",
						 "100011011110001111010010",
						 "100011011110010011000010",
						 "100011011110010110110010",
						 "100011011110011010100010",
						 "100011011101100010010010",
						 "100011011101100110000010",
						 "100011011101101001110010",
						 "100011011101101101100010",
						 "100011011101110001010010",
						 "100011011101110101000010",
						 "100011011101111000110010",
						 "100011011101111100100010",
						 "100011011110000000010010",
						 "100011011110000100000010",
						 "100011011110000111110010",
						 "100011011110001011100010",
						 "100011011110001111010010",
						 "100011011110010011000010",
						 "100011011110010110110010",
						 "100011011110011010100010",
						 "100011011101100010010010",
						 "100011011101100110000001",
						 "100011011101101001110000",
						 "100011011101101101011111",
						 "100011011101110001001110",
						 "100011011101110100111101",
						 "100011011101111000101100",
						 "100011011101111100011011",
						 "100011011110000000001010",
						 "100011011110000011111001",
						 "100011011110000111101000",
						 "100011011110001011010111",
						 "100011011110001111000110",
						 "100011011110010010110101",
						 "100011011110010110100100",
						 "100011011110011010010011",
						 "100011100000000101010000",
						 "100011100000001000111111",
						 "100011100000001100101110",
						 "100011100000010000011101",
						 "100011100000010100001100",
						 "100011100000010111111011",
						 "100011100000011011101010",
						 "100011100000011111011001",
						 "100011100000100011001000",
						 "100011100000100110110111",
						 "100011100000101010100110",
						 "100011100000101110010101",
						 "100011100000110010000100",
						 "100011100000110101110011",
						 "100011100000111001100010",
						 "100011100000111101010001",
						 "100011100000000101010000",
						 "100011100000001000111111",
						 "100011100000001100101110",
						 "100011100000010000011101",
						 "100011100000010100001100",
						 "100011100000010111111011",
						 "100011100000011011101010",
						 "100011100000011111011001",
						 "100011100000100011001000",
						 "100011100000100110110111",
						 "100011100000101010100110",
						 "100011100000101110010101",
						 "100011100000110010000100",
						 "100011100000110101110011",
						 "100011100000111001100010",
						 "100011100000111101010001",
						 "100011100000000101010000",
						 "100011100000001000111111",
						 "100011100000001100101110",
						 "100011100000010000011101",
						 "100011100000010100001100",
						 "100011100000010111111011",
						 "100011100000011011101010",
						 "100011100000011111011001",
						 "100011100000100011001000",
						 "100011100000100110110111",
						 "100011100000101010100110",
						 "100011100000101110010101",
						 "100011100000110010000100",
						 "100011100000110101110011",
						 "100011100000111001100010",
						 "100011100000111101010001",
						 "100011100010101000001110",
						 "100011100010101011111101",
						 "100011100010101111101100",
						 "100011100010110011011011",
						 "100011100010110111001010",
						 "100011100010111010111001",
						 "100011100010111110101000",
						 "100011100011000010010111",
						 "100011100011000110000110",
						 "100011100011001001110101",
						 "100011100011001101100100",
						 "100011100011010001010011",
						 "100011100011010101000010",
						 "100011100011011000110001",
						 "100011100011011100100000",
						 "100011100011100000001111",
						 "100011100010101000001110",
						 "100011100010101011111101",
						 "100011100010101111101100",
						 "100011100010110011011011",
						 "100011100010110111001010",
						 "100011100010111010111001",
						 "100011100010111110101000",
						 "100011100011000010010111",
						 "100011100011000110000110",
						 "100011100011001001110101",
						 "100011100011001101100100",
						 "100011100011010001010011",
						 "100011100011010101000010",
						 "100011100011011000110001",
						 "100011100011011100100000",
						 "100011100011100000001111",
						 "100011100101001011001100",
						 "100011100101001110111011",
						 "100011100101010010101010",
						 "100011100101010110011001",
						 "100011100101011010001000",
						 "100011100101011101110111",
						 "100011100101100001100110",
						 "100011100101100101010101",
						 "100011100101101001000100",
						 "100011100101101100110011",
						 "100011100101110000100010",
						 "100011100101110100010001",
						 "100011100101111000000000",
						 "100011100101111011101111",
						 "100011100101111111011110",
						 "100011100110000011001101",
						 "100011100101001011001100",
						 "100011100101001110111011",
						 "100011100101010010101010",
						 "100011100101010110011001",
						 "100011100101011010001000",
						 "100011100101011101110111",
						 "100011100101100001100110",
						 "100011100101100101010101",
						 "100011100101101001000100",
						 "100011100101101100110011",
						 "100011100101110000100010",
						 "100011100101110100010001",
						 "100011100101111000000000",
						 "100011100101111011101111",
						 "100011100101111111011110",
						 "100011100110000011001101",
						 "100011100101001011001100",
						 "100011100101001110111010",
						 "100011100101010010101000",
						 "100011100101010110010110",
						 "100011100101011010000100",
						 "100011100101011101110010",
						 "100011100101100001100000",
						 "100011100101100101001110",
						 "100011100101101000111100",
						 "100011100101101100101010",
						 "100011100101110000011000",
						 "100011100101110100000110",
						 "100011100101110111110100",
						 "100011100101111011100010",
						 "100011100101111111010000",
						 "100011100110000010111110",
						 "100011100111101110001010",
						 "100011100111110001111000",
						 "100011100111110101100110",
						 "100011100111111001010100",
						 "100011100111111101000010",
						 "100011101000000000110000",
						 "100011101000000100011110",
						 "100011101000001000001100",
						 "100011101000001011111010",
						 "100011101000001111101000",
						 "100011101000010011010110",
						 "100011101000010111000100",
						 "100011101000011010110010",
						 "100011101000011110100000",
						 "100011101000100010001110",
						 "100011101000100101111100",
						 "100011100111101110001010",
						 "100011100111110001111000",
						 "100011100111110101100110",
						 "100011100111111001010100",
						 "100011100111111101000010",
						 "100011101000000000110000",
						 "100011101000000100011110",
						 "100011101000001000001100",
						 "100011101000001011111010",
						 "100011101000001111101000",
						 "100011101000010011010110",
						 "100011101000010111000100",
						 "100011101000011010110010",
						 "100011101000011110100000",
						 "100011101000100010001110",
						 "100011101000100101111100",
						 "100011100111101110001010",
						 "100011100111110001111000",
						 "100011100111110101100110",
						 "100011100111111001010100",
						 "100011100111111101000010",
						 "100011101000000000110000",
						 "100011101000000100011110",
						 "100011101000001000001100",
						 "100011101000001011111010",
						 "100011101000001111101000",
						 "100011101000010011010110",
						 "100011101000010111000100",
						 "100011101000011010110010",
						 "100011101000011110100000",
						 "100011101000100010001110",
						 "100011101000100101111100",
						 "100011101010010001001000",
						 "100011101010010100110110",
						 "100011101010011000100100",
						 "100011101010011100010010",
						 "100011101010100000000000",
						 "100011101010100011101110",
						 "100011101010100111011100",
						 "100011101010101011001010",
						 "100011101010101110111000",
						 "100011101010110010100110",
						 "100011101010110110010100",
						 "100011101010111010000010",
						 "100011101010111101110000",
						 "100011101011000001011110",
						 "100011101011000101001100",
						 "100011101011001000111010",
						 "100011101010010001001000",
						 "100011101010010100110110",
						 "100011101010011000100100",
						 "100011101010011100010010",
						 "100011101010100000000000",
						 "100011101010100011101110",
						 "100011101010100111011100",
						 "100011101010101011001010",
						 "100011101010101110111000",
						 "100011101010110010100110",
						 "100011101010110110010100",
						 "100011101010111010000010",
						 "100011101010111101110000",
						 "100011101011000001011110",
						 "100011101011000101001100",
						 "100011101011001000111010",
						 "100011101100110100000110",
						 "100011101100110111110100",
						 "100011101100111011100010",
						 "100011101100111111010000",
						 "100011101101000010111110",
						 "100011101101000110101100",
						 "100011101101001010011010",
						 "100011101101001110001000",
						 "100011101101010001110110",
						 "100011101101010101100100",
						 "100011101101011001010010",
						 "100011101101011101000000",
						 "100011101101100000101110",
						 "100011101101100100011100",
						 "100011101101101000001010",
						 "100011101101101011111000",
						 "100011101100110100000110",
						 "100011101100110111110011",
						 "100011101100111011100000",
						 "100011101100111111001101",
						 "100011101101000010111010",
						 "100011101101000110100111",
						 "100011101101001010010100",
						 "100011101101001110000001",
						 "100011101101010001101110",
						 "100011101101010101011011",
						 "100011101101011001001000",
						 "100011101101011100110101",
						 "100011101101100000100010",
						 "100011101101100100001111",
						 "100011101101100111111100",
						 "100011101101101011101001",
						 "100011101100110100000110",
						 "100011101100110111110011",
						 "100011101100111011100000",
						 "100011101100111111001101",
						 "100011101101000010111010",
						 "100011101101000110100111",
						 "100011101101001010010100",
						 "100011101101001110000001",
						 "100011101101010001101110",
						 "100011101101010101011011",
						 "100011101101011001001000",
						 "100011101101011100110101",
						 "100011101101100000100010",
						 "100011101101100100001111",
						 "100011101101100111111100",
						 "100011101101101011101001",
						 "100011101111010111000100",
						 "100011101111011010110001",
						 "100011101111011110011110",
						 "100011101111100010001011",
						 "100011101111100101111000",
						 "100011101111101001100101",
						 "100011101111101101010010",
						 "100011101111110000111111",
						 "100011101111110100101100",
						 "100011101111111000011001",
						 "100011101111111100000110",
						 "100011101111111111110011",
						 "100011110000000011100000",
						 "100011110000000111001101",
						 "100011110000001010111010",
						 "100011110000001110100111",
						 "100011101111010111000100",
						 "100011101111011010110001",
						 "100011101111011110011110",
						 "100011101111100010001011",
						 "100011101111100101111000",
						 "100011101111101001100101",
						 "100011101111101101010010",
						 "100011101111110000111111",
						 "100011101111110100101100",
						 "100011101111111000011001",
						 "100011101111111100000110",
						 "100011101111111111110011",
						 "100011110000000011100000",
						 "100011110000000111001101",
						 "100011110000001010111010",
						 "100011110000001110100111",
						 "100011101111010111000100",
						 "100011101111011010110001",
						 "100011101111011110011110",
						 "100011101111100010001011",
						 "100011101111100101111000",
						 "100011101111101001100101",
						 "100011101111101101010010",
						 "100011101111110000111111",
						 "100011101111110100101100",
						 "100011101111111000011001",
						 "100011101111111100000110",
						 "100011101111111111110011",
						 "100011110000000011100000",
						 "100011110000000111001101",
						 "100011110000001010111010",
						 "100011110000001110100111",
						 "100011110001111010000010",
						 "100011110001111101101111",
						 "100011110010000001011100",
						 "100011110010000101001001",
						 "100011110010001000110110",
						 "100011110010001100100011",
						 "100011110010010000010000",
						 "100011110010010011111101",
						 "100011110010010111101010",
						 "100011110010011011010111",
						 "100011110010011111000100",
						 "100011110010100010110001",
						 "100011110010100110011110",
						 "100011110010101010001011",
						 "100011110010101101111000",
						 "100011110010110001100101",
						 "100011110001111010000010",
						 "100011110001111101101111",
						 "100011110010000001011100",
						 "100011110010000101001001",
						 "100011110010001000110110",
						 "100011110010001100100011",
						 "100011110010010000010000",
						 "100011110010010011111101",
						 "100011110010010111101010",
						 "100011110010011011010111",
						 "100011110010011111000100",
						 "100011110010100010110001",
						 "100011110010100110011110",
						 "100011110010101010001011",
						 "100011110010101101111000",
						 "100011110010110001100101",
						 "100011110001111010000010",
						 "100011110001111101101110",
						 "100011110010000001011010",
						 "100011110010000101000110",
						 "100011110010001000110010",
						 "100011110010001100011110",
						 "100011110010010000001010",
						 "100011110010010011110110",
						 "100011110010010111100010",
						 "100011110010011011001110",
						 "100011110010011110111010",
						 "100011110010100010100110",
						 "100011110010100110010010",
						 "100011110010101001111110",
						 "100011110010101101101010",
						 "100011110010110001010110",
						 "100011110100011101000000",
						 "100011110100100000101100",
						 "100011110100100100011000",
						 "100011110100101000000100",
						 "100011110100101011110000",
						 "100011110100101111011100",
						 "100011110100110011001000",
						 "100011110100110110110100",
						 "100011110100111010100000",
						 "100011110100111110001100",
						 "100011110101000001111000",
						 "100011110101000101100100",
						 "100011110101001001010000",
						 "100011110101001100111100",
						 "100011110101010000101000",
						 "100011110101010100010100",
						 "100011110100011101000000",
						 "100011110100100000101100",
						 "100011110100100100011000",
						 "100011110100101000000100",
						 "100011110100101011110000",
						 "100011110100101111011100",
						 "100011110100110011001000",
						 "100011110100110110110100",
						 "100011110100111010100000",
						 "100011110100111110001100",
						 "100011110101000001111000",
						 "100011110101000101100100",
						 "100011110101001001010000",
						 "100011110101001100111100",
						 "100011110101010000101000",
						 "100011110101010100010100",
						 "100011110110111111111110",
						 "100011110111000011101010",
						 "100011110111000111010110",
						 "100011110111001011000010",
						 "100011110111001110101110",
						 "100011110111010010011010",
						 "100011110111010110000110",
						 "100011110111011001110010",
						 "100011110111011101011110",
						 "100011110111100001001010",
						 "100011110111100100110110",
						 "100011110111101000100010",
						 "100011110111101100001110",
						 "100011110111101111111010",
						 "100011110111110011100110",
						 "100011110111110111010010",
						 "100011110110111111111110",
						 "100011110111000011101010",
						 "100011110111000111010110",
						 "100011110111001011000010",
						 "100011110111001110101110",
						 "100011110111010010011010",
						 "100011110111010110000110",
						 "100011110111011001110010",
						 "100011110111011101011110",
						 "100011110111100001001010",
						 "100011110111100100110110",
						 "100011110111101000100010",
						 "100011110111101100001110",
						 "100011110111101111111010",
						 "100011110111110011100110",
						 "100011110111110111010010",
						 "100011110110111111111110",
						 "100011110111000011101010",
						 "100011110111000111010110",
						 "100011110111001011000010",
						 "100011110111001110101110",
						 "100011110111010010011010",
						 "100011110111010110000110",
						 "100011110111011001110010",
						 "100011110111011101011110",
						 "100011110111100001001010",
						 "100011110111100100110110",
						 "100011110111101000100010",
						 "100011110111101100001110",
						 "100011110111101111111010",
						 "100011110111110011100110",
						 "100011110111110111010010",
						 "100011111001100010111100",
						 "100011111001100110101000",
						 "100011111001101010010100",
						 "100011111001101110000000",
						 "100011111001110001101100",
						 "100011111001110101011000",
						 "100011111001111001000100",
						 "100011111001111100110000",
						 "100011111010000000011100",
						 "100011111010000100001000",
						 "100011111010000111110100",
						 "100011111010001011100000",
						 "100011111010001111001100",
						 "100011111010010010111000",
						 "100011111010010110100100",
						 "100011111010011010010000",
						 "100011111001100010111100",
						 "100011111001100110100111",
						 "100011111001101010010010",
						 "100011111001101101111101",
						 "100011111001110001101000",
						 "100011111001110101010011",
						 "100011111001111000111110",
						 "100011111001111100101001",
						 "100011111010000000010100",
						 "100011111010000011111111",
						 "100011111010000111101010",
						 "100011111010001011010101",
						 "100011111010001111000000",
						 "100011111010010010101011",
						 "100011111010010110010110",
						 "100011111010011010000001",
						 "100011111001100010111100",
						 "100011111001100110100111",
						 "100011111001101010010010",
						 "100011111001101101111101",
						 "100011111001110001101000",
						 "100011111001110101010011",
						 "100011111001111000111110",
						 "100011111001111100101001",
						 "100011111010000000010100",
						 "100011111010000011111111",
						 "100011111010000111101010",
						 "100011111010001011010101",
						 "100011111010001111000000",
						 "100011111010010010101011",
						 "100011111010010110010110",
						 "100011111010011010000001",
						 "100011111100000101111010",
						 "100011111100001001100101",
						 "100011111100001101010000",
						 "100011111100010000111011",
						 "100011111100010100100110",
						 "100011111100011000010001",
						 "100011111100011011111100",
						 "100011111100011111100111",
						 "100011111100100011010010",
						 "100011111100100110111101",
						 "100011111100101010101000",
						 "100011111100101110010011",
						 "100011111100110001111110",
						 "100011111100110101101001",
						 "100011111100111001010100",
						 "100011111100111100111111",
						 "100011111100000101111010",
						 "100011111100001001100101",
						 "100011111100001101010000",
						 "100011111100010000111011",
						 "100011111100010100100110",
						 "100011111100011000010001",
						 "100011111100011011111100",
						 "100011111100011111100111",
						 "100011111100100011010010",
						 "100011111100100110111101",
						 "100011111100101010101000",
						 "100011111100101110010011",
						 "100011111100110001111110",
						 "100011111100110101101001",
						 "100011111100111001010100",
						 "100011111100111100111111",
						 "100011111100000101111010",
						 "100011111100001001100101",
						 "100011111100001101010000",
						 "100011111100010000111011",
						 "100011111100010100100110",
						 "100011111100011000010001",
						 "100011111100011011111100",
						 "100011111100011111100111",
						 "100011111100100011010010",
						 "100011111100100110111101",
						 "100011111100101010101000",
						 "100011111100101110010011",
						 "100011111100110001111110",
						 "100011111100110101101001",
						 "100011111100111001010100",
						 "100011111100111100111111",
						 "100011111110101000111000",
						 "100011111110101100100011",
						 "100011111110110000001110",
						 "100011111110110011111001",
						 "100011111110110111100100",
						 "100011111110111011001111",
						 "100011111110111110111010",
						 "100011111111000010100101",
						 "100011111111000110010000",
						 "100011111111001001111011",
						 "100011111111001101100110",
						 "100011111111010001010001",
						 "100011111111010100111100",
						 "100011111111011000100111",
						 "100011111111011100010010",
						 "100011111111011111111101",
						 "100011111110101000111000",
						 "100011111110101100100010",
						 "100011111110110000001100",
						 "100011111110110011110110",
						 "100011111110110111100000",
						 "100011111110111011001010",
						 "100011111110111110110100",
						 "100011111111000010011110",
						 "100011111111000110001000",
						 "100011111111001001110010",
						 "100011111111001101011100",
						 "100011111111010001000110",
						 "100011111111010100110000",
						 "100011111111011000011010",
						 "100011111111011100000100",
						 "100011111111011111101110",
						 "100011111110101000111000",
						 "100011111110101100100010",
						 "100011111110110000001100",
						 "100011111110110011110110",
						 "100011111110110111100000",
						 "100011111110111011001010",
						 "100011111110111110110100",
						 "100011111111000010011110",
						 "100011111111000110001000",
						 "100011111111001001110010",
						 "100011111111001101011100",
						 "100011111111010001000110",
						 "100011111111010100110000",
						 "100011111111011000011010",
						 "100011111111011100000100",
						 "100011111111011111101110",
						 "100100000001001011110110",
						 "100100000001001111100000",
						 "100100000001010011001010",
						 "100100000001010110110100",
						 "100100000001011010011110",
						 "100100000001011110001000",
						 "100100000001100001110010",
						 "100100000001100101011100",
						 "100100000001101001000110",
						 "100100000001101100110000",
						 "100100000001110000011010",
						 "100100000001110100000100",
						 "100100000001110111101110",
						 "100100000001111011011000",
						 "100100000001111111000010",
						 "100100000010000010101100",
						 "100100000001001011110110",
						 "100100000001001111100000",
						 "100100000001010011001010",
						 "100100000001010110110100",
						 "100100000001011010011110",
						 "100100000001011110001000",
						 "100100000001100001110010",
						 "100100000001100101011100",
						 "100100000001101001000110",
						 "100100000001101100110000",
						 "100100000001110000011010",
						 "100100000001110100000100",
						 "100100000001110111101110",
						 "100100000001111011011000",
						 "100100000001111111000010",
						 "100100000010000010101100",
						 "100100000011101110110100",
						 "100100000011110010011110",
						 "100100000011110110001000",
						 "100100000011111001110010",
						 "100100000011111101011100",
						 "100100000100000001000110",
						 "100100000100000100110000",
						 "100100000100001000011010",
						 "100100000100001100000100",
						 "100100000100001111101110",
						 "100100000100010011011000",
						 "100100000100010111000010",
						 "100100000100011010101100",
						 "100100000100011110010110",
						 "100100000100100010000000",
						 "100100000100100101101010",
						 "100100000011101110110100",
						 "100100000011110010011110",
						 "100100000011110110001000",
						 "100100000011111001110010",
						 "100100000011111101011100",
						 "100100000100000001000110",
						 "100100000100000100110000",
						 "100100000100001000011010",
						 "100100000100001100000100",
						 "100100000100001111101110",
						 "100100000100010011011000",
						 "100100000100010111000010",
						 "100100000100011010101100",
						 "100100000100011110010110",
						 "100100000100100010000000",
						 "100100000100100101101010",
						 "100100000011101110110100",
						 "100100000011110010011110",
						 "100100000011110110001000",
						 "100100000011111001110010",
						 "100100000011111101011100",
						 "100100000100000001000110",
						 "100100000100000100110000",
						 "100100000100001000011010",
						 "100100000100001100000100",
						 "100100000100001111101110",
						 "100100000100010011011000",
						 "100100000100010111000010",
						 "100100000100011010101100",
						 "100100000100011110010110",
						 "100100000100100010000000",
						 "100100000100100101101010",
						 "100100000110010001110010",
						 "100100000110010101011011",
						 "100100000110011001000100",
						 "100100000110011100101101",
						 "100100000110100000010110",
						 "100100000110100011111111",
						 "100100000110100111101000",
						 "100100000110101011010001",
						 "100100000110101110111010",
						 "100100000110110010100011",
						 "100100000110110110001100",
						 "100100000110111001110101",
						 "100100000110111101011110",
						 "100100000111000001000111",
						 "100100000111000100110000",
						 "100100000111001000011001",
						 "100100000110010001110010",
						 "100100000110010101011011",
						 "100100000110011001000100",
						 "100100000110011100101101",
						 "100100000110100000010110",
						 "100100000110100011111111",
						 "100100000110100111101000",
						 "100100000110101011010001",
						 "100100000110101110111010",
						 "100100000110110010100011",
						 "100100000110110110001100",
						 "100100000110111001110101",
						 "100100000110111101011110",
						 "100100000111000001000111",
						 "100100000111000100110000",
						 "100100000111001000011001",
						 "100100000110010001110010",
						 "100100000110010101011011",
						 "100100000110011001000100",
						 "100100000110011100101101",
						 "100100000110100000010110",
						 "100100000110100011111111",
						 "100100000110100111101000",
						 "100100000110101011010001",
						 "100100000110101110111010",
						 "100100000110110010100011",
						 "100100000110110110001100",
						 "100100000110111001110101",
						 "100100000110111101011110",
						 "100100000111000001000111",
						 "100100000111000100110000",
						 "100100000111001000011001",
						 "100100001000110100110000",
						 "100100001000111000011001",
						 "100100001000111100000010",
						 "100100001000111111101011",
						 "100100001001000011010100",
						 "100100001001000110111101",
						 "100100001001001010100110",
						 "100100001001001110001111",
						 "100100001001010001111000",
						 "100100001001010101100001",
						 "100100001001011001001010",
						 "100100001001011100110011",
						 "100100001001100000011100",
						 "100100001001100100000101",
						 "100100001001100111101110",
						 "100100001001101011010111",
						 "100100001000110100110000",
						 "100100001000111000011001",
						 "100100001000111100000010",
						 "100100001000111111101011",
						 "100100001001000011010100",
						 "100100001001000110111101",
						 "100100001001001010100110",
						 "100100001001001110001111",
						 "100100001001010001111000",
						 "100100001001010101100001",
						 "100100001001011001001010",
						 "100100001001011100110011",
						 "100100001001100000011100",
						 "100100001001100100000101",
						 "100100001001100111101110",
						 "100100001001101011010111",
						 "100100001000110100110000",
						 "100100001000111000011001",
						 "100100001000111100000010",
						 "100100001000111111101011",
						 "100100001001000011010100",
						 "100100001001000110111101",
						 "100100001001001010100110",
						 "100100001001001110001111",
						 "100100001001010001111000",
						 "100100001001010101100001",
						 "100100001001011001001010",
						 "100100001001011100110011",
						 "100100001001100000011100",
						 "100100001001100100000101",
						 "100100001001100111101110",
						 "100100001001101011010111",
						 "100100001011010111101110",
						 "100100001011011011010110",
						 "100100001011011110111110",
						 "100100001011100010100110",
						 "100100001011100110001110",
						 "100100001011101001110110",
						 "100100001011101101011110",
						 "100100001011110001000110",
						 "100100001011110100101110",
						 "100100001011111000010110",
						 "100100001011111011111110",
						 "100100001011111111100110",
						 "100100001100000011001110",
						 "100100001100000110110110",
						 "100100001100001010011110",
						 "100100001100001110000110",
						 "100100001011010111101110",
						 "100100001011011011010110",
						 "100100001011011110111110",
						 "100100001011100010100110",
						 "100100001011100110001110",
						 "100100001011101001110110",
						 "100100001011101101011110",
						 "100100001011110001000110",
						 "100100001011110100101110",
						 "100100001011111000010110",
						 "100100001011111011111110",
						 "100100001011111111100110",
						 "100100001100000011001110",
						 "100100001100000110110110",
						 "100100001100001010011110",
						 "100100001100001110000110",
						 "100100001011010111101110",
						 "100100001011011011010110",
						 "100100001011011110111110",
						 "100100001011100010100110",
						 "100100001011100110001110",
						 "100100001011101001110110",
						 "100100001011101101011110",
						 "100100001011110001000110",
						 "100100001011110100101110",
						 "100100001011111000010110",
						 "100100001011111011111110",
						 "100100001011111111100110",
						 "100100001100000011001110",
						 "100100001100000110110110",
						 "100100001100001010011110",
						 "100100001100001110000110",
						 "100100001101111010101100",
						 "100100001101111110010100",
						 "100100001110000001111100",
						 "100100001110000101100100",
						 "100100001110001001001100",
						 "100100001110001100110100",
						 "100100001110010000011100",
						 "100100001110010100000100",
						 "100100001110010111101100",
						 "100100001110011011010100",
						 "100100001110011110111100",
						 "100100001110100010100100",
						 "100100001110100110001100",
						 "100100001110101001110100",
						 "100100001110101101011100",
						 "100100001110110001000100",
						 "100100001101111010101100",
						 "100100001101111110010100",
						 "100100001110000001111100",
						 "100100001110000101100100",
						 "100100001110001001001100",
						 "100100001110001100110100",
						 "100100001110010000011100",
						 "100100001110010100000100",
						 "100100001110010111101100",
						 "100100001110011011010100",
						 "100100001110011110111100",
						 "100100001110100010100100",
						 "100100001110100110001100",
						 "100100001110101001110100",
						 "100100001110101101011100",
						 "100100001110110001000100",
						 "100100010000011101101010",
						 "100100010000100001010010",
						 "100100010000100100111010",
						 "100100010000101000100010",
						 "100100010000101100001010",
						 "100100010000101111110010",
						 "100100010000110011011010",
						 "100100010000110111000010",
						 "100100010000111010101010",
						 "100100010000111110010010",
						 "100100010001000001111010",
						 "100100010001000101100010",
						 "100100010001001001001010",
						 "100100010001001100110010",
						 "100100010001010000011010",
						 "100100010001010100000010",
						 "100100010000011101101010",
						 "100100010000100001010001",
						 "100100010000100100111000",
						 "100100010000101000011111",
						 "100100010000101100000110",
						 "100100010000101111101101",
						 "100100010000110011010100",
						 "100100010000110110111011",
						 "100100010000111010100010",
						 "100100010000111110001001",
						 "100100010001000001110000",
						 "100100010001000101010111",
						 "100100010001001000111110",
						 "100100010001001100100101",
						 "100100010001010000001100",
						 "100100010001010011110011",
						 "100100010000011101101010",
						 "100100010000100001010001",
						 "100100010000100100111000",
						 "100100010000101000011111",
						 "100100010000101100000110",
						 "100100010000101111101101",
						 "100100010000110011010100",
						 "100100010000110110111011",
						 "100100010000111010100010",
						 "100100010000111110001001",
						 "100100010001000001110000",
						 "100100010001000101010111",
						 "100100010001001000111110",
						 "100100010001001100100101",
						 "100100010001010000001100",
						 "100100010001010011110011",
						 "100100010011000000101000",
						 "100100010011000100001111",
						 "100100010011000111110110",
						 "100100010011001011011101",
						 "100100010011001111000100",
						 "100100010011010010101011",
						 "100100010011010110010010",
						 "100100010011011001111001",
						 "100100010011011101100000",
						 "100100010011100001000111",
						 "100100010011100100101110",
						 "100100010011101000010101",
						 "100100010011101011111100",
						 "100100010011101111100011",
						 "100100010011110011001010",
						 "100100010011110110110001",
						 "100100010011000000101000",
						 "100100010011000100001111",
						 "100100010011000111110110",
						 "100100010011001011011101",
						 "100100010011001111000100",
						 "100100010011010010101011",
						 "100100010011010110010010",
						 "100100010011011001111001",
						 "100100010011011101100000",
						 "100100010011100001000111",
						 "100100010011100100101110",
						 "100100010011101000010101",
						 "100100010011101011111100",
						 "100100010011101111100011",
						 "100100010011110011001010",
						 "100100010011110110110001",
						 "100100010011000000101000",
						 "100100010011000100001111",
						 "100100010011000111110110",
						 "100100010011001011011101",
						 "100100010011001111000100",
						 "100100010011010010101011",
						 "100100010011010110010010",
						 "100100010011011001111001",
						 "100100010011011101100000",
						 "100100010011100001000111",
						 "100100010011100100101110",
						 "100100010011101000010101",
						 "100100010011101011111100",
						 "100100010011101111100011",
						 "100100010011110011001010",
						 "100100010011110110110001",
						 "100100010101100011100110",
						 "100100010101100111001101",
						 "100100010101101010110100",
						 "100100010101101110011011",
						 "100100010101110010000010",
						 "100100010101110101101001",
						 "100100010101111001010000",
						 "100100010101111100110111",
						 "100100010110000000011110",
						 "100100010110000100000101",
						 "100100010110000111101100",
						 "100100010110001011010011",
						 "100100010110001110111010",
						 "100100010110010010100001",
						 "100100010110010110001000",
						 "100100010110011001101111",
						 "100100010101100011100110",
						 "100100010101100111001100",
						 "100100010101101010110010",
						 "100100010101101110011000",
						 "100100010101110001111110",
						 "100100010101110101100100",
						 "100100010101111001001010",
						 "100100010101111100110000",
						 "100100010110000000010110",
						 "100100010110000011111100",
						 "100100010110000111100010",
						 "100100010110001011001000",
						 "100100010110001110101110",
						 "100100010110010010010100",
						 "100100010110010101111010",
						 "100100010110011001100000",
						 "100100010101100011100110",
						 "100100010101100111001100",
						 "100100010101101010110010",
						 "100100010101101110011000",
						 "100100010101110001111110",
						 "100100010101110101100100",
						 "100100010101111001001010",
						 "100100010101111100110000",
						 "100100010110000000010110",
						 "100100010110000011111100",
						 "100100010110000111100010",
						 "100100010110001011001000",
						 "100100010110001110101110",
						 "100100010110010010010100",
						 "100100010110010101111010",
						 "100100010110011001100000",
						 "100100011000000110100100",
						 "100100011000001010001010",
						 "100100011000001101110000",
						 "100100011000010001010110",
						 "100100011000010100111100",
						 "100100011000011000100010",
						 "100100011000011100001000",
						 "100100011000011111101110",
						 "100100011000100011010100",
						 "100100011000100110111010",
						 "100100011000101010100000",
						 "100100011000101110000110",
						 "100100011000110001101100",
						 "100100011000110101010010",
						 "100100011000111000111000",
						 "100100011000111100011110",
						 "100100011000000110100100",
						 "100100011000001010001010",
						 "100100011000001101110000",
						 "100100011000010001010110",
						 "100100011000010100111100",
						 "100100011000011000100010",
						 "100100011000011100001000",
						 "100100011000011111101110",
						 "100100011000100011010100",
						 "100100011000100110111010",
						 "100100011000101010100000",
						 "100100011000101110000110",
						 "100100011000110001101100",
						 "100100011000110101010010",
						 "100100011000111000111000",
						 "100100011000111100011110",
						 "100100011000000110100100",
						 "100100011000001010001010",
						 "100100011000001101110000",
						 "100100011000010001010110",
						 "100100011000010100111100",
						 "100100011000011000100010",
						 "100100011000011100001000",
						 "100100011000011111101110",
						 "100100011000100011010100",
						 "100100011000100110111010",
						 "100100011000101010100000",
						 "100100011000101110000110",
						 "100100011000110001101100",
						 "100100011000110101010010",
						 "100100011000111000111000",
						 "100100011000111100011110",
						 "100100011010101001100010",
						 "100100011010101101001000",
						 "100100011010110000101110",
						 "100100011010110100010100",
						 "100100011010110111111010",
						 "100100011010111011100000",
						 "100100011010111111000110",
						 "100100011011000010101100",
						 "100100011011000110010010",
						 "100100011011001001111000",
						 "100100011011001101011110",
						 "100100011011010001000100",
						 "100100011011010100101010",
						 "100100011011011000010000",
						 "100100011011011011110110",
						 "100100011011011111011100",
						 "100100011010101001100010",
						 "100100011010101101000111",
						 "100100011010110000101100",
						 "100100011010110100010001",
						 "100100011010110111110110",
						 "100100011010111011011011",
						 "100100011010111111000000",
						 "100100011011000010100101",
						 "100100011011000110001010",
						 "100100011011001001101111",
						 "100100011011001101010100",
						 "100100011011010000111001",
						 "100100011011010100011110",
						 "100100011011011000000011",
						 "100100011011011011101000",
						 "100100011011011111001101",
						 "100100011010101001100010",
						 "100100011010101101000111",
						 "100100011010110000101100",
						 "100100011010110100010001",
						 "100100011010110111110110",
						 "100100011010111011011011",
						 "100100011010111111000000",
						 "100100011011000010100101",
						 "100100011011000110001010",
						 "100100011011001001101111",
						 "100100011011001101010100",
						 "100100011011010000111001",
						 "100100011011010100011110",
						 "100100011011011000000011",
						 "100100011011011011101000",
						 "100100011011011111001101",
						 "100100011101001100100000",
						 "100100011101010000000101",
						 "100100011101010011101010",
						 "100100011101010111001111",
						 "100100011101011010110100",
						 "100100011101011110011001",
						 "100100011101100001111110",
						 "100100011101100101100011",
						 "100100011101101001001000",
						 "100100011101101100101101",
						 "100100011101110000010010",
						 "100100011101110011110111",
						 "100100011101110111011100",
						 "100100011101111011000001",
						 "100100011101111110100110",
						 "100100011110000010001011",
						 "100100011101001100100000",
						 "100100011101010000000101",
						 "100100011101010011101010",
						 "100100011101010111001111",
						 "100100011101011010110100",
						 "100100011101011110011001",
						 "100100011101100001111110",
						 "100100011101100101100011",
						 "100100011101101001001000",
						 "100100011101101100101101",
						 "100100011101110000010010",
						 "100100011101110011110111",
						 "100100011101110111011100",
						 "100100011101111011000001",
						 "100100011101111110100110",
						 "100100011110000010001011",
						 "100100011111101111011110",
						 "100100011111110011000011",
						 "100100011111110110101000",
						 "100100011111111010001101",
						 "100100011111111101110010",
						 "100100100000000001010111",
						 "100100100000000100111100",
						 "100100100000001000100001",
						 "100100100000001100000110",
						 "100100100000001111101011",
						 "100100100000010011010000",
						 "100100100000010110110101",
						 "100100100000011010011010",
						 "100100100000011101111111",
						 "100100100000100001100100",
						 "100100100000100101001001",
						 "100100011111101111011110",
						 "100100011111110011000011",
						 "100100011111110110101000",
						 "100100011111111010001101",
						 "100100011111111101110010",
						 "100100100000000001010111",
						 "100100100000000100111100",
						 "100100100000001000100001",
						 "100100100000001100000110",
						 "100100100000001111101011",
						 "100100100000010011010000",
						 "100100100000010110110101",
						 "100100100000011010011010",
						 "100100100000011101111111",
						 "100100100000100001100100",
						 "100100100000100101001001",
						 "100100011111101111011110",
						 "100100011111110011000010",
						 "100100011111110110100110",
						 "100100011111111010001010",
						 "100100011111111101101110",
						 "100100100000000001010010",
						 "100100100000000100110110",
						 "100100100000001000011010",
						 "100100100000001011111110",
						 "100100100000001111100010",
						 "100100100000010011000110",
						 "100100100000010110101010",
						 "100100100000011010001110",
						 "100100100000011101110010",
						 "100100100000100001010110",
						 "100100100000100100111010",
						 "100100100010010010011100",
						 "100100100010010110000000",
						 "100100100010011001100100",
						 "100100100010011101001000",
						 "100100100010100000101100",
						 "100100100010100100010000",
						 "100100100010100111110100",
						 "100100100010101011011000",
						 "100100100010101110111100",
						 "100100100010110010100000",
						 "100100100010110110000100",
						 "100100100010111001101000",
						 "100100100010111101001100",
						 "100100100011000000110000",
						 "100100100011000100010100",
						 "100100100011000111111000",
						 "100100100010010010011100",
						 "100100100010010110000000",
						 "100100100010011001100100",
						 "100100100010011101001000",
						 "100100100010100000101100",
						 "100100100010100100010000",
						 "100100100010100111110100",
						 "100100100010101011011000",
						 "100100100010101110111100",
						 "100100100010110010100000",
						 "100100100010110110000100",
						 "100100100010111001101000",
						 "100100100010111101001100",
						 "100100100011000000110000",
						 "100100100011000100010100",
						 "100100100011000111111000",
						 "100100100010010010011100",
						 "100100100010010110000000",
						 "100100100010011001100100",
						 "100100100010011101001000",
						 "100100100010100000101100",
						 "100100100010100100010000",
						 "100100100010100111110100",
						 "100100100010101011011000",
						 "100100100010101110111100",
						 "100100100010110010100000",
						 "100100100010110110000100",
						 "100100100010111001101000",
						 "100100100010111101001100",
						 "100100100011000000110000",
						 "100100100011000100010100",
						 "100100100011000111111000",
						 "100100100100110101011010",
						 "100100100100111000111110",
						 "100100100100111100100010",
						 "100100100101000000000110",
						 "100100100101000011101010",
						 "100100100101000111001110",
						 "100100100101001010110010",
						 "100100100101001110010110",
						 "100100100101010001111010",
						 "100100100101010101011110",
						 "100100100101011001000010",
						 "100100100101011100100110",
						 "100100100101100000001010",
						 "100100100101100011101110",
						 "100100100101100111010010",
						 "100100100101101010110110",
						 "100100100100110101011010",
						 "100100100100111000111110",
						 "100100100100111100100010",
						 "100100100101000000000110",
						 "100100100101000011101010",
						 "100100100101000111001110",
						 "100100100101001010110010",
						 "100100100101001110010110",
						 "100100100101010001111010",
						 "100100100101010101011110",
						 "100100100101011001000010",
						 "100100100101011100100110",
						 "100100100101100000001010",
						 "100100100101100011101110",
						 "100100100101100111010010",
						 "100100100101101010110110",
						 "100100100100110101011010",
						 "100100100100111000111101",
						 "100100100100111100100000",
						 "100100100101000000000011",
						 "100100100101000011100110",
						 "100100100101000111001001",
						 "100100100101001010101100",
						 "100100100101001110001111",
						 "100100100101010001110010",
						 "100100100101010101010101",
						 "100100100101011000111000",
						 "100100100101011100011011",
						 "100100100101011111111110",
						 "100100100101100011100001",
						 "100100100101100111000100",
						 "100100100101101010100111",
						 "100100100111011000011000",
						 "100100100111011011111011",
						 "100100100111011111011110",
						 "100100100111100011000001",
						 "100100100111100110100100",
						 "100100100111101010000111",
						 "100100100111101101101010",
						 "100100100111110001001101",
						 "100100100111110100110000",
						 "100100100111111000010011",
						 "100100100111111011110110",
						 "100100100111111111011001",
						 "100100101000000010111100",
						 "100100101000000110011111",
						 "100100101000001010000010",
						 "100100101000001101100101",
						 "100100100111011000011000",
						 "100100100111011011111011",
						 "100100100111011111011110",
						 "100100100111100011000001",
						 "100100100111100110100100",
						 "100100100111101010000111",
						 "100100100111101101101010",
						 "100100100111110001001101",
						 "100100100111110100110000",
						 "100100100111111000010011",
						 "100100100111111011110110",
						 "100100100111111111011001",
						 "100100101000000010111100",
						 "100100101000000110011111",
						 "100100101000001010000010",
						 "100100101000001101100101",
						 "100100100111011000011000",
						 "100100100111011011111011",
						 "100100100111011111011110",
						 "100100100111100011000001",
						 "100100100111100110100100",
						 "100100100111101010000111",
						 "100100100111101101101010",
						 "100100100111110001001101",
						 "100100100111110100110000",
						 "100100100111111000010011",
						 "100100100111111011110110",
						 "100100100111111111011001",
						 "100100101000000010111100",
						 "100100101000000110011111",
						 "100100101000001010000010",
						 "100100101000001101100101",
						 "100100101001111011010110",
						 "100100101001111110111001",
						 "100100101010000010011100",
						 "100100101010000101111111",
						 "100100101010001001100010",
						 "100100101010001101000101",
						 "100100101010010000101000",
						 "100100101010010100001011",
						 "100100101010010111101110",
						 "100100101010011011010001",
						 "100100101010011110110100",
						 "100100101010100010010111",
						 "100100101010100101111010",
						 "100100101010101001011101",
						 "100100101010101101000000",
						 "100100101010110000100011",
						 "100100101001111011010110",
						 "100100101001111110111000",
						 "100100101010000010011010",
						 "100100101010000101111100",
						 "100100101010001001011110",
						 "100100101010001101000000",
						 "100100101010010000100010",
						 "100100101010010100000100",
						 "100100101010010111100110",
						 "100100101010011011001000",
						 "100100101010011110101010",
						 "100100101010100010001100",
						 "100100101010100101101110",
						 "100100101010101001010000",
						 "100100101010101100110010",
						 "100100101010110000010100",
						 "100100101001111011010110",
						 "100100101001111110111000",
						 "100100101010000010011010",
						 "100100101010000101111100",
						 "100100101010001001011110",
						 "100100101010001101000000",
						 "100100101010010000100010",
						 "100100101010010100000100",
						 "100100101010010111100110",
						 "100100101010011011001000",
						 "100100101010011110101010",
						 "100100101010100010001100",
						 "100100101010100101101110",
						 "100100101010101001010000",
						 "100100101010101100110010",
						 "100100101010110000010100",
						 "100100101100011110010100",
						 "100100101100100001110110",
						 "100100101100100101011000",
						 "100100101100101000111010",
						 "100100101100101100011100",
						 "100100101100101111111110",
						 "100100101100110011100000",
						 "100100101100110111000010",
						 "100100101100111010100100",
						 "100100101100111110000110",
						 "100100101101000001101000",
						 "100100101101000101001010",
						 "100100101101001000101100",
						 "100100101101001100001110",
						 "100100101101001111110000",
						 "100100101101010011010010",
						 "100100101100011110010100",
						 "100100101100100001110110",
						 "100100101100100101011000",
						 "100100101100101000111010",
						 "100100101100101100011100",
						 "100100101100101111111110",
						 "100100101100110011100000",
						 "100100101100110111000010",
						 "100100101100111010100100",
						 "100100101100111110000110",
						 "100100101101000001101000",
						 "100100101101000101001010",
						 "100100101101001000101100",
						 "100100101101001100001110",
						 "100100101101001111110000",
						 "100100101101010011010010",
						 "100100101100011110010100",
						 "100100101100100001110110",
						 "100100101100100101011000",
						 "100100101100101000111010",
						 "100100101100101100011100",
						 "100100101100101111111110",
						 "100100101100110011100000",
						 "100100101100110111000010",
						 "100100101100111010100100",
						 "100100101100111110000110",
						 "100100101101000001101000",
						 "100100101101000101001010",
						 "100100101101001000101100",
						 "100100101101001100001110",
						 "100100101101001111110000",
						 "100100101101010011010010",
						 "100100101111000001010010",
						 "100100101111000100110100",
						 "100100101111001000010110",
						 "100100101111001011111000",
						 "100100101111001111011010",
						 "100100101111010010111100",
						 "100100101111010110011110",
						 "100100101111011010000000",
						 "100100101111011101100010",
						 "100100101111100001000100",
						 "100100101111100100100110",
						 "100100101111101000001000",
						 "100100101111101011101010",
						 "100100101111101111001100",
						 "100100101111110010101110",
						 "100100101111110110010000",
						 "100100101111000001010010",
						 "100100101111000100110011",
						 "100100101111001000010100",
						 "100100101111001011110101",
						 "100100101111001111010110",
						 "100100101111010010110111",
						 "100100101111010110011000",
						 "100100101111011001111001",
						 "100100101111011101011010",
						 "100100101111100000111011",
						 "100100101111100100011100",
						 "100100101111100111111101",
						 "100100101111101011011110",
						 "100100101111101110111111",
						 "100100101111110010100000",
						 "100100101111110110000001",
						 "100100110001100100010000",
						 "100100110001100111110001",
						 "100100110001101011010010",
						 "100100110001101110110011",
						 "100100110001110010010100",
						 "100100110001110101110101",
						 "100100110001111001010110",
						 "100100110001111100110111",
						 "100100110010000000011000",
						 "100100110010000011111001",
						 "100100110010000111011010",
						 "100100110010001010111011",
						 "100100110010001110011100",
						 "100100110010010001111101",
						 "100100110010010101011110",
						 "100100110010011000111111",
						 "100100110001100100010000",
						 "100100110001100111110001",
						 "100100110001101011010010",
						 "100100110001101110110011",
						 "100100110001110010010100",
						 "100100110001110101110101",
						 "100100110001111001010110",
						 "100100110001111100110111",
						 "100100110010000000011000",
						 "100100110010000011111001",
						 "100100110010000111011010",
						 "100100110010001010111011",
						 "100100110010001110011100",
						 "100100110010010001111101",
						 "100100110010010101011110",
						 "100100110010011000111111",
						 "100100110001100100010000",
						 "100100110001100111110001",
						 "100100110001101011010010",
						 "100100110001101110110011",
						 "100100110001110010010100",
						 "100100110001110101110101",
						 "100100110001111001010110",
						 "100100110001111100110111",
						 "100100110010000000011000",
						 "100100110010000011111001",
						 "100100110010000111011010",
						 "100100110010001010111011",
						 "100100110010001110011100",
						 "100100110010010001111101",
						 "100100110010010101011110",
						 "100100110010011000111111",
						 "100100110100000111001110",
						 "100100110100001010101111",
						 "100100110100001110010000",
						 "100100110100010001110001",
						 "100100110100010101010010",
						 "100100110100011000110011",
						 "100100110100011100010100",
						 "100100110100011111110101",
						 "100100110100100011010110",
						 "100100110100100110110111",
						 "100100110100101010011000",
						 "100100110100101101111001",
						 "100100110100110001011010",
						 "100100110100110100111011",
						 "100100110100111000011100",
						 "100100110100111011111101",
						 "100100110100000111001110",
						 "100100110100001010101110",
						 "100100110100001110001110",
						 "100100110100010001101110",
						 "100100110100010101001110",
						 "100100110100011000101110",
						 "100100110100011100001110",
						 "100100110100011111101110",
						 "100100110100100011001110",
						 "100100110100100110101110",
						 "100100110100101010001110",
						 "100100110100101101101110",
						 "100100110100110001001110",
						 "100100110100110100101110",
						 "100100110100111000001110",
						 "100100110100111011101110",
						 "100100110100000111001110",
						 "100100110100001010101110",
						 "100100110100001110001110",
						 "100100110100010001101110",
						 "100100110100010101001110",
						 "100100110100011000101110",
						 "100100110100011100001110",
						 "100100110100011111101110",
						 "100100110100100011001110",
						 "100100110100100110101110",
						 "100100110100101010001110",
						 "100100110100101101101110",
						 "100100110100110001001110",
						 "100100110100110100101110",
						 "100100110100111000001110",
						 "100100110100111011101110",
						 "100100110110101010001100",
						 "100100110110101101101100",
						 "100100110110110001001100",
						 "100100110110110100101100",
						 "100100110110111000001100",
						 "100100110110111011101100",
						 "100100110110111111001100",
						 "100100110111000010101100",
						 "100100110111000110001100",
						 "100100110111001001101100",
						 "100100110111001101001100",
						 "100100110111010000101100",
						 "100100110111010100001100",
						 "100100110111010111101100",
						 "100100110111011011001100",
						 "100100110111011110101100",
						 "100100110110101010001100",
						 "100100110110101101101100",
						 "100100110110110001001100",
						 "100100110110110100101100",
						 "100100110110111000001100",
						 "100100110110111011101100",
						 "100100110110111111001100",
						 "100100110111000010101100",
						 "100100110111000110001100",
						 "100100110111001001101100",
						 "100100110111001101001100",
						 "100100110111010000101100",
						 "100100110111010100001100",
						 "100100110111010111101100",
						 "100100110111011011001100",
						 "100100110111011110101100",
						 "100100110110101010001100",
						 "100100110110101101101100",
						 "100100110110110001001100",
						 "100100110110110100101100",
						 "100100110110111000001100",
						 "100100110110111011101100",
						 "100100110110111111001100",
						 "100100110111000010101100",
						 "100100110111000110001100",
						 "100100110111001001101100",
						 "100100110111001101001100",
						 "100100110111010000101100",
						 "100100110111010100001100",
						 "100100110111010111101100",
						 "100100110111011011001100",
						 "100100110111011110101100",
						 "100100111001001101001010",
						 "100100111001010000101001",
						 "100100111001010100001000",
						 "100100111001010111100111",
						 "100100111001011011000110",
						 "100100111001011110100101",
						 "100100111001100010000100",
						 "100100111001100101100011",
						 "100100111001101001000010",
						 "100100111001101100100001",
						 "100100111001110000000000",
						 "100100111001110011011111",
						 "100100111001110110111110",
						 "100100111001111010011101",
						 "100100111001111101111100",
						 "100100111010000001011011",
						 "100100111001001101001010",
						 "100100111001010000101001",
						 "100100111001010100001000",
						 "100100111001010111100111",
						 "100100111001011011000110",
						 "100100111001011110100101",
						 "100100111001100010000100",
						 "100100111001100101100011",
						 "100100111001101001000010",
						 "100100111001101100100001",
						 "100100111001110000000000",
						 "100100111001110011011111",
						 "100100111001110110111110",
						 "100100111001111010011101",
						 "100100111001111101111100",
						 "100100111010000001011011",
						 "100100111001001101001010",
						 "100100111001010000101001",
						 "100100111001010100001000",
						 "100100111001010111100111",
						 "100100111001011011000110",
						 "100100111001011110100101",
						 "100100111001100010000100",
						 "100100111001100101100011",
						 "100100111001101001000010",
						 "100100111001101100100001",
						 "100100111001110000000000",
						 "100100111001110011011111",
						 "100100111001110110111110",
						 "100100111001111010011101",
						 "100100111001111101111100",
						 "100100111010000001011011",
						 "100100111011110000001000",
						 "100100111011110011100111",
						 "100100111011110111000110",
						 "100100111011111010100101",
						 "100100111011111110000100",
						 "100100111100000001100011",
						 "100100111100000101000010",
						 "100100111100001000100001",
						 "100100111100001100000000",
						 "100100111100001111011111",
						 "100100111100010010111110",
						 "100100111100010110011101",
						 "100100111100011001111100",
						 "100100111100011101011011",
						 "100100111100100000111010",
						 "100100111100100100011001",
						 "100100111011110000001000",
						 "100100111011110011100111",
						 "100100111011110111000110",
						 "100100111011111010100101",
						 "100100111011111110000100",
						 "100100111100000001100011",
						 "100100111100000101000010",
						 "100100111100001000100001",
						 "100100111100001100000000",
						 "100100111100001111011111",
						 "100100111100010010111110",
						 "100100111100010110011101",
						 "100100111100011001111100",
						 "100100111100011101011011",
						 "100100111100100000111010",
						 "100100111100100100011001",
						 "100100111011110000001000",
						 "100100111011110011100111",
						 "100100111011110111000110",
						 "100100111011111010100101",
						 "100100111011111110000100",
						 "100100111100000001100011",
						 "100100111100000101000010",
						 "100100111100001000100001",
						 "100100111100001100000000",
						 "100100111100001111011111",
						 "100100111100010010111110",
						 "100100111100010110011101",
						 "100100111100011001111100",
						 "100100111100011101011011",
						 "100100111100100000111010",
						 "100100111100100100011001",
						 "100100111110010011000110",
						 "100100111110010110100100",
						 "100100111110011010000010",
						 "100100111110011101100000",
						 "100100111110100000111110",
						 "100100111110100100011100",
						 "100100111110100111111010",
						 "100100111110101011011000",
						 "100100111110101110110110",
						 "100100111110110010010100",
						 "100100111110110101110010",
						 "100100111110111001010000",
						 "100100111110111100101110",
						 "100100111111000000001100",
						 "100100111111000011101010",
						 "100100111111000111001000",
						 "100100111110010011000110",
						 "100100111110010110100100",
						 "100100111110011010000010",
						 "100100111110011101100000",
						 "100100111110100000111110",
						 "100100111110100100011100",
						 "100100111110100111111010",
						 "100100111110101011011000",
						 "100100111110101110110110",
						 "100100111110110010010100",
						 "100100111110110101110010",
						 "100100111110111001010000",
						 "100100111110111100101110",
						 "100100111111000000001100",
						 "100100111111000011101010",
						 "100100111111000111001000",
						 "100100111110010011000110",
						 "100100111110010110100100",
						 "100100111110011010000010",
						 "100100111110011101100000",
						 "100100111110100000111110",
						 "100100111110100100011100",
						 "100100111110100111111010",
						 "100100111110101011011000",
						 "100100111110101110110110",
						 "100100111110110010010100",
						 "100100111110110101110010",
						 "100100111110111001010000",
						 "100100111110111100101110",
						 "100100111111000000001100",
						 "100100111111000011101010",
						 "100100111111000111001000",
						 "100101000000110110000100",
						 "100101000000111001100010",
						 "100101000000111101000000",
						 "100101000001000000011110",
						 "100101000001000011111100",
						 "100101000001000111011010",
						 "100101000001001010111000",
						 "100101000001001110010110",
						 "100101000001010001110100",
						 "100101000001010101010010",
						 "100101000001011000110000",
						 "100101000001011100001110",
						 "100101000001011111101100",
						 "100101000001100011001010",
						 "100101000001100110101000",
						 "100101000001101010000110",
						 "100101000000110110000100",
						 "100101000000111001100010",
						 "100101000000111101000000",
						 "100101000001000000011110",
						 "100101000001000011111100",
						 "100101000001000111011010",
						 "100101000001001010111000",
						 "100101000001001110010110",
						 "100101000001010001110100",
						 "100101000001010101010010",
						 "100101000001011000110000",
						 "100101000001011100001110",
						 "100101000001011111101100",
						 "100101000001100011001010",
						 "100101000001100110101000",
						 "100101000001101010000110",
						 "100101000000110110000100",
						 "100101000000111001100001",
						 "100101000000111100111110",
						 "100101000001000000011011",
						 "100101000001000011111000",
						 "100101000001000111010101",
						 "100101000001001010110010",
						 "100101000001001110001111",
						 "100101000001010001101100",
						 "100101000001010101001001",
						 "100101000001011000100110",
						 "100101000001011100000011",
						 "100101000001011111100000",
						 "100101000001100010111101",
						 "100101000001100110011010",
						 "100101000001101001110111",
						 "100101000011011001000010",
						 "100101000011011100011111",
						 "100101000011011111111100",
						 "100101000011100011011001",
						 "100101000011100110110110",
						 "100101000011101010010011",
						 "100101000011101101110000",
						 "100101000011110001001101",
						 "100101000011110100101010",
						 "100101000011111000000111",
						 "100101000011111011100100",
						 "100101000011111111000001",
						 "100101000100000010011110",
						 "100101000100000101111011",
						 "100101000100001001011000",
						 "100101000100001100110101",
						 "100101000011011001000010",
						 "100101000011011100011111",
						 "100101000011011111111100",
						 "100101000011100011011001",
						 "100101000011100110110110",
						 "100101000011101010010011",
						 "100101000011101101110000",
						 "100101000011110001001101",
						 "100101000011110100101010",
						 "100101000011111000000111",
						 "100101000011111011100100",
						 "100101000011111111000001",
						 "100101000100000010011110",
						 "100101000100000101111011",
						 "100101000100001001011000",
						 "100101000100001100110101",
						 "100101000011011001000010",
						 "100101000011011100011111",
						 "100101000011011111111100",
						 "100101000011100011011001",
						 "100101000011100110110110",
						 "100101000011101010010011",
						 "100101000011101101110000",
						 "100101000011110001001101",
						 "100101000011110100101010",
						 "100101000011111000000111",
						 "100101000011111011100100",
						 "100101000011111111000001",
						 "100101000100000010011110",
						 "100101000100000101111011",
						 "100101000100001001011000",
						 "100101000100001100110101",
						 "100101000101111100000000",
						 "100101000101111111011101",
						 "100101000110000010111010",
						 "100101000110000110010111",
						 "100101000110001001110100",
						 "100101000110001101010001",
						 "100101000110010000101110",
						 "100101000110010100001011",
						 "100101000110010111101000",
						 "100101000110011011000101",
						 "100101000110011110100010",
						 "100101000110100001111111",
						 "100101000110100101011100",
						 "100101000110101000111001",
						 "100101000110101100010110",
						 "100101000110101111110011",
						 "100101000101111100000000",
						 "100101000101111111011100",
						 "100101000110000010111000",
						 "100101000110000110010100",
						 "100101000110001001110000",
						 "100101000110001101001100",
						 "100101000110010000101000",
						 "100101000110010100000100",
						 "100101000110010111100000",
						 "100101000110011010111100",
						 "100101000110011110011000",
						 "100101000110100001110100",
						 "100101000110100101010000",
						 "100101000110101000101100",
						 "100101000110101100001000",
						 "100101000110101111100100",
						 "100101000101111100000000",
						 "100101000101111111011100",
						 "100101000110000010111000",
						 "100101000110000110010100",
						 "100101000110001001110000",
						 "100101000110001101001100",
						 "100101000110010000101000",
						 "100101000110010100000100",
						 "100101000110010111100000",
						 "100101000110011010111100",
						 "100101000110011110011000",
						 "100101000110100001110100",
						 "100101000110100101010000",
						 "100101000110101000101100",
						 "100101000110101100001000",
						 "100101000110101111100100",
						 "100101001000011110111110",
						 "100101001000100010011010",
						 "100101001000100101110110",
						 "100101001000101001010010",
						 "100101001000101100101110",
						 "100101001000110000001010",
						 "100101001000110011100110",
						 "100101001000110111000010",
						 "100101001000111010011110",
						 "100101001000111101111010",
						 "100101001001000001010110",
						 "100101001001000100110010",
						 "100101001001001000001110",
						 "100101001001001011101010",
						 "100101001001001111000110",
						 "100101001001010010100010",
						 "100101001000011110111110",
						 "100101001000100010011010",
						 "100101001000100101110110",
						 "100101001000101001010010",
						 "100101001000101100101110",
						 "100101001000110000001010",
						 "100101001000110011100110",
						 "100101001000110111000010",
						 "100101001000111010011110",
						 "100101001000111101111010",
						 "100101001001000001010110",
						 "100101001001000100110010",
						 "100101001001001000001110",
						 "100101001001001011101010",
						 "100101001001001111000110",
						 "100101001001010010100010",
						 "100101001000011110111110",
						 "100101001000100010011010",
						 "100101001000100101110110",
						 "100101001000101001010010",
						 "100101001000101100101110",
						 "100101001000110000001010",
						 "100101001000110011100110",
						 "100101001000110111000010",
						 "100101001000111010011110",
						 "100101001000111101111010",
						 "100101001001000001010110",
						 "100101001001000100110010",
						 "100101001001001000001110",
						 "100101001001001011101010",
						 "100101001001001111000110",
						 "100101001001010010100010",
						 "100101001011000001111100",
						 "100101001011000101010111",
						 "100101001011001000110010",
						 "100101001011001100001101",
						 "100101001011001111101000",
						 "100101001011010011000011",
						 "100101001011010110011110",
						 "100101001011011001111001",
						 "100101001011011101010100",
						 "100101001011100000101111",
						 "100101001011100100001010",
						 "100101001011100111100101",
						 "100101001011101011000000",
						 "100101001011101110011011",
						 "100101001011110001110110",
						 "100101001011110101010001",
						 "100101001011000001111100",
						 "100101001011000101010111",
						 "100101001011001000110010",
						 "100101001011001100001101",
						 "100101001011001111101000",
						 "100101001011010011000011",
						 "100101001011010110011110",
						 "100101001011011001111001",
						 "100101001011011101010100",
						 "100101001011100000101111",
						 "100101001011100100001010",
						 "100101001011100111100101",
						 "100101001011101011000000",
						 "100101001011101110011011",
						 "100101001011110001110110",
						 "100101001011110101010001",
						 "100101001011000001111100",
						 "100101001011000101010111",
						 "100101001011001000110010",
						 "100101001011001100001101",
						 "100101001011001111101000",
						 "100101001011010011000011",
						 "100101001011010110011110",
						 "100101001011011001111001",
						 "100101001011011101010100",
						 "100101001011100000101111",
						 "100101001011100100001010",
						 "100101001011100111100101",
						 "100101001011101011000000",
						 "100101001011101110011011",
						 "100101001011110001110110",
						 "100101001011110101010001",
						 "100101001101100100111010",
						 "100101001101101000010101",
						 "100101001101101011110000",
						 "100101001101101111001011",
						 "100101001101110010100110",
						 "100101001101110110000001",
						 "100101001101111001011100",
						 "100101001101111100110111",
						 "100101001110000000010010",
						 "100101001110000011101101",
						 "100101001110000111001000",
						 "100101001110001010100011",
						 "100101001110001101111110",
						 "100101001110010001011001",
						 "100101001110010100110100",
						 "100101001110011000001111",
						 "100101001101100100111010",
						 "100101001101101000010101",
						 "100101001101101011110000",
						 "100101001101101111001011",
						 "100101001101110010100110",
						 "100101001101110110000001",
						 "100101001101111001011100",
						 "100101001101111100110111",
						 "100101001110000000010010",
						 "100101001110000011101101",
						 "100101001110000111001000",
						 "100101001110001010100011",
						 "100101001110001101111110",
						 "100101001110010001011001",
						 "100101001110010100110100",
						 "100101001110011000001111",
						 "100101001101100100111010",
						 "100101001101101000010100",
						 "100101001101101011101110",
						 "100101001101101111001000",
						 "100101001101110010100010",
						 "100101001101110101111100",
						 "100101001101111001010110",
						 "100101001101111100110000",
						 "100101001110000000001010",
						 "100101001110000011100100",
						 "100101001110000110111110",
						 "100101001110001010011000",
						 "100101001110001101110010",
						 "100101001110010001001100",
						 "100101001110010100100110",
						 "100101001110011000000000",
						 "100101010000000111111000",
						 "100101010000001011010010",
						 "100101010000001110101100",
						 "100101010000010010000110",
						 "100101010000010101100000",
						 "100101010000011000111010",
						 "100101010000011100010100",
						 "100101010000011111101110",
						 "100101010000100011001000",
						 "100101010000100110100010",
						 "100101010000101001111100",
						 "100101010000101101010110",
						 "100101010000110000110000",
						 "100101010000110100001010",
						 "100101010000110111100100",
						 "100101010000111010111110",
						 "100101010000000111111000",
						 "100101010000001011010010",
						 "100101010000001110101100",
						 "100101010000010010000110",
						 "100101010000010101100000",
						 "100101010000011000111010",
						 "100101010000011100010100",
						 "100101010000011111101110",
						 "100101010000100011001000",
						 "100101010000100110100010",
						 "100101010000101001111100",
						 "100101010000101101010110",
						 "100101010000110000110000",
						 "100101010000110100001010",
						 "100101010000110111100100",
						 "100101010000111010111110",
						 "100101010000000111111000",
						 "100101010000001011010010",
						 "100101010000001110101100",
						 "100101010000010010000110",
						 "100101010000010101100000",
						 "100101010000011000111010",
						 "100101010000011100010100",
						 "100101010000011111101110",
						 "100101010000100011001000",
						 "100101010000100110100010",
						 "100101010000101001111100",
						 "100101010000101101010110",
						 "100101010000110000110000",
						 "100101010000110100001010",
						 "100101010000110111100100",
						 "100101010000111010111110",
						 "100101010010101010110110",
						 "100101010010101110010000",
						 "100101010010110001101010",
						 "100101010010110101000100",
						 "100101010010111000011110",
						 "100101010010111011111000",
						 "100101010010111111010010",
						 "100101010011000010101100",
						 "100101010011000110000110",
						 "100101010011001001100000",
						 "100101010011001100111010",
						 "100101010011010000010100",
						 "100101010011010011101110",
						 "100101010011010111001000",
						 "100101010011011010100010",
						 "100101010011011101111100",
						 "100101010010101010110110",
						 "100101010010101110001111",
						 "100101010010110001101000",
						 "100101010010110101000001",
						 "100101010010111000011010",
						 "100101010010111011110011",
						 "100101010010111111001100",
						 "100101010011000010100101",
						 "100101010011000101111110",
						 "100101010011001001010111",
						 "100101010011001100110000",
						 "100101010011010000001001",
						 "100101010011010011100010",
						 "100101010011010110111011",
						 "100101010011011010010100",
						 "100101010011011101101101",
						 "100101010010101010110110",
						 "100101010010101110001111",
						 "100101010010110001101000",
						 "100101010010110101000001",
						 "100101010010111000011010",
						 "100101010010111011110011",
						 "100101010010111111001100",
						 "100101010011000010100101",
						 "100101010011000101111110",
						 "100101010011001001010111",
						 "100101010011001100110000",
						 "100101010011010000001001",
						 "100101010011010011100010",
						 "100101010011010110111011",
						 "100101010011011010010100",
						 "100101010011011101101101",
						 "100101010101001101110100",
						 "100101010101010001001101",
						 "100101010101010100100110",
						 "100101010101010111111111",
						 "100101010101011011011000",
						 "100101010101011110110001",
						 "100101010101100010001010",
						 "100101010101100101100011",
						 "100101010101101000111100",
						 "100101010101101100010101",
						 "100101010101101111101110",
						 "100101010101110011000111",
						 "100101010101110110100000",
						 "100101010101111001111001",
						 "100101010101111101010010",
						 "100101010110000000101011",
						 "100101010101001101110100",
						 "100101010101010001001101",
						 "100101010101010100100110",
						 "100101010101010111111111",
						 "100101010101011011011000",
						 "100101010101011110110001",
						 "100101010101100010001010",
						 "100101010101100101100011",
						 "100101010101101000111100",
						 "100101010101101100010101",
						 "100101010101101111101110",
						 "100101010101110011000111",
						 "100101010101110110100000",
						 "100101010101111001111001",
						 "100101010101111101010010",
						 "100101010110000000101011",
						 "100101010101001101110100",
						 "100101010101010001001101",
						 "100101010101010100100110",
						 "100101010101010111111111",
						 "100101010101011011011000",
						 "100101010101011110110001",
						 "100101010101100010001010",
						 "100101010101100101100011",
						 "100101010101101000111100",
						 "100101010101101100010101",
						 "100101010101101111101110",
						 "100101010101110011000111",
						 "100101010101110110100000",
						 "100101010101111001111001",
						 "100101010101111101010010",
						 "100101010110000000101011",
						 "100101010111110000110010",
						 "100101010111110100001010",
						 "100101010111110111100010",
						 "100101010111111010111010",
						 "100101010111111110010010",
						 "100101011000000001101010",
						 "100101011000000101000010",
						 "100101011000001000011010",
						 "100101011000001011110010",
						 "100101011000001111001010",
						 "100101011000010010100010",
						 "100101011000010101111010",
						 "100101011000011001010010",
						 "100101011000011100101010",
						 "100101011000100000000010",
						 "100101011000100011011010",
						 "100101010111110000110010",
						 "100101010111110100001010",
						 "100101010111110111100010",
						 "100101010111111010111010",
						 "100101010111111110010010",
						 "100101011000000001101010",
						 "100101011000000101000010",
						 "100101011000001000011010",
						 "100101011000001011110010",
						 "100101011000001111001010",
						 "100101011000010010100010",
						 "100101011000010101111010",
						 "100101011000011001010010",
						 "100101011000011100101010",
						 "100101011000100000000010",
						 "100101011000100011011010",
						 "100101010111110000110010",
						 "100101010111110100001010",
						 "100101010111110111100010",
						 "100101010111111010111010",
						 "100101010111111110010010",
						 "100101011000000001101010",
						 "100101011000000101000010",
						 "100101011000001000011010",
						 "100101011000001011110010",
						 "100101011000001111001010",
						 "100101011000010010100010",
						 "100101011000010101111010",
						 "100101011000011001010010",
						 "100101011000011100101010",
						 "100101011000100000000010",
						 "100101011000100011011010",
						 "100101011010010011110000",
						 "100101011010010111001000",
						 "100101011010011010100000",
						 "100101011010011101111000",
						 "100101011010100001010000",
						 "100101011010100100101000",
						 "100101011010101000000000",
						 "100101011010101011011000",
						 "100101011010101110110000",
						 "100101011010110010001000",
						 "100101011010110101100000",
						 "100101011010111000111000",
						 "100101011010111100010000",
						 "100101011010111111101000",
						 "100101011011000011000000",
						 "100101011011000110011000",
						 "100101011010010011110000",
						 "100101011010010111001000",
						 "100101011010011010100000",
						 "100101011010011101111000",
						 "100101011010100001010000",
						 "100101011010100100101000",
						 "100101011010101000000000",
						 "100101011010101011011000",
						 "100101011010101110110000",
						 "100101011010110010001000",
						 "100101011010110101100000",
						 "100101011010111000111000",
						 "100101011010111100010000",
						 "100101011010111111101000",
						 "100101011011000011000000",
						 "100101011011000110011000",
						 "100101011010010011110000",
						 "100101011010010111000111",
						 "100101011010011010011110",
						 "100101011010011101110101",
						 "100101011010100001001100",
						 "100101011010100100100011",
						 "100101011010100111111010",
						 "100101011010101011010001",
						 "100101011010101110101000",
						 "100101011010110001111111",
						 "100101011010110101010110",
						 "100101011010111000101101",
						 "100101011010111100000100",
						 "100101011010111111011011",
						 "100101011011000010110010",
						 "100101011011000110001001",
						 "100101011100110110101110",
						 "100101011100111010000101",
						 "100101011100111101011100",
						 "100101011101000000110011",
						 "100101011101000100001010",
						 "100101011101000111100001",
						 "100101011101001010111000",
						 "100101011101001110001111",
						 "100101011101010001100110",
						 "100101011101010100111101",
						 "100101011101011000010100",
						 "100101011101011011101011",
						 "100101011101011111000010",
						 "100101011101100010011001",
						 "100101011101100101110000",
						 "100101011101101001000111",
						 "100101011100110110101110",
						 "100101011100111010000101",
						 "100101011100111101011100",
						 "100101011101000000110011",
						 "100101011101000100001010",
						 "100101011101000111100001",
						 "100101011101001010111000",
						 "100101011101001110001111",
						 "100101011101010001100110",
						 "100101011101010100111101",
						 "100101011101011000010100",
						 "100101011101011011101011",
						 "100101011101011111000010",
						 "100101011101100010011001",
						 "100101011101100101110000",
						 "100101011101101001000111",
						 "100101011100110110101110",
						 "100101011100111010000101",
						 "100101011100111101011100",
						 "100101011101000000110011",
						 "100101011101000100001010",
						 "100101011101000111100001",
						 "100101011101001010111000",
						 "100101011101001110001111",
						 "100101011101010001100110",
						 "100101011101010100111101",
						 "100101011101011000010100",
						 "100101011101011011101011",
						 "100101011101011111000010",
						 "100101011101100010011001",
						 "100101011101100101110000",
						 "100101011101101001000111",
						 "100101011111011001101100",
						 "100101011111011101000010",
						 "100101011111100000011000",
						 "100101011111100011101110",
						 "100101011111100111000100",
						 "100101011111101010011010",
						 "100101011111101101110000",
						 "100101011111110001000110",
						 "100101011111110100011100",
						 "100101011111110111110010",
						 "100101011111111011001000",
						 "100101011111111110011110",
						 "100101100000000001110100",
						 "100101100000000101001010",
						 "100101100000001000100000",
						 "100101100000001011110110",
						 "100101011111011001101100",
						 "100101011111011101000010",
						 "100101011111100000011000",
						 "100101011111100011101110",
						 "100101011111100111000100",
						 "100101011111101010011010",
						 "100101011111101101110000",
						 "100101011111110001000110",
						 "100101011111110100011100",
						 "100101011111110111110010",
						 "100101011111111011001000",
						 "100101011111111110011110",
						 "100101100000000001110100",
						 "100101100000000101001010",
						 "100101100000001000100000",
						 "100101100000001011110110",
						 "100101011111011001101100",
						 "100101011111011101000010",
						 "100101011111100000011000",
						 "100101011111100011101110",
						 "100101011111100111000100",
						 "100101011111101010011010",
						 "100101011111101101110000",
						 "100101011111110001000110",
						 "100101011111110100011100",
						 "100101011111110111110010",
						 "100101011111111011001000",
						 "100101011111111110011110",
						 "100101100000000001110100",
						 "100101100000000101001010",
						 "100101100000001000100000",
						 "100101100000001011110110",
						 "100101100001111100101010",
						 "100101100010000000000000",
						 "100101100010000011010110",
						 "100101100010000110101100",
						 "100101100010001010000010",
						 "100101100010001101011000",
						 "100101100010010000101110",
						 "100101100010010100000100",
						 "100101100010010111011010",
						 "100101100010011010110000",
						 "100101100010011110000110",
						 "100101100010100001011100",
						 "100101100010100100110010",
						 "100101100010101000001000",
						 "100101100010101011011110",
						 "100101100010101110110100",
						 "100101100001111100101010",
						 "100101100010000000000000",
						 "100101100010000011010110",
						 "100101100010000110101100",
						 "100101100010001010000010",
						 "100101100010001101011000",
						 "100101100010010000101110",
						 "100101100010010100000100",
						 "100101100010010111011010",
						 "100101100010011010110000",
						 "100101100010011110000110",
						 "100101100010100001011100",
						 "100101100010100100110010",
						 "100101100010101000001000",
						 "100101100010101011011110",
						 "100101100010101110110100",
						 "100101100001111100101010",
						 "100101100001111111111111",
						 "100101100010000011010100",
						 "100101100010000110101001",
						 "100101100010001001111110",
						 "100101100010001101010011",
						 "100101100010010000101000",
						 "100101100010010011111101",
						 "100101100010010111010010",
						 "100101100010011010100111",
						 "100101100010011101111100",
						 "100101100010100001010001",
						 "100101100010100100100110",
						 "100101100010100111111011",
						 "100101100010101011010000",
						 "100101100010101110100101",
						 "100101100100011111101000",
						 "100101100100100010111101",
						 "100101100100100110010010",
						 "100101100100101001100111",
						 "100101100100101100111100",
						 "100101100100110000010001",
						 "100101100100110011100110",
						 "100101100100110110111011",
						 "100101100100111010010000",
						 "100101100100111101100101",
						 "100101100101000000111010",
						 "100101100101000100001111",
						 "100101100101000111100100",
						 "100101100101001010111001",
						 "100101100101001110001110",
						 "100101100101010001100011",
						 "100101100100011111101000",
						 "100101100100100010111101",
						 "100101100100100110010010",
						 "100101100100101001100111",
						 "100101100100101100111100",
						 "100101100100110000010001",
						 "100101100100110011100110",
						 "100101100100110110111011",
						 "100101100100111010010000",
						 "100101100100111101100101",
						 "100101100101000000111010",
						 "100101100101000100001111",
						 "100101100101000111100100",
						 "100101100101001010111001",
						 "100101100101001110001110",
						 "100101100101010001100011",
						 "100101100100011111101000",
						 "100101100100100010111101",
						 "100101100100100110010010",
						 "100101100100101001100111",
						 "100101100100101100111100",
						 "100101100100110000010001",
						 "100101100100110011100110",
						 "100101100100110110111011",
						 "100101100100111010010000",
						 "100101100100111101100101",
						 "100101100101000000111010",
						 "100101100101000100001111",
						 "100101100101000111100100",
						 "100101100101001010111001",
						 "100101100101001110001110",
						 "100101100101010001100011",
						 "100101100111000010100110",
						 "100101100111000101111011",
						 "100101100111001001010000",
						 "100101100111001100100101",
						 "100101100111001111111010",
						 "100101100111010011001111",
						 "100101100111010110100100",
						 "100101100111011001111001",
						 "100101100111011101001110",
						 "100101100111100000100011",
						 "100101100111100011111000",
						 "100101100111100111001101",
						 "100101100111101010100010",
						 "100101100111101101110111",
						 "100101100111110001001100",
						 "100101100111110100100001",
						 "100101100111000010100110",
						 "100101100111000101111010",
						 "100101100111001001001110",
						 "100101100111001100100010",
						 "100101100111001111110110",
						 "100101100111010011001010",
						 "100101100111010110011110",
						 "100101100111011001110010",
						 "100101100111011101000110",
						 "100101100111100000011010",
						 "100101100111100011101110",
						 "100101100111100111000010",
						 "100101100111101010010110",
						 "100101100111101101101010",
						 "100101100111110000111110",
						 "100101100111110100010010",
						 "100101100111000010100110",
						 "100101100111000101111010",
						 "100101100111001001001110",
						 "100101100111001100100010",
						 "100101100111001111110110",
						 "100101100111010011001010",
						 "100101100111010110011110",
						 "100101100111011001110010",
						 "100101100111011101000110",
						 "100101100111100000011010",
						 "100101100111100011101110",
						 "100101100111100111000010",
						 "100101100111101010010110",
						 "100101100111101101101010",
						 "100101100111110000111110",
						 "100101100111110100010010",
						 "100101101001100101100100",
						 "100101101001101000111000",
						 "100101101001101100001100",
						 "100101101001101111100000",
						 "100101101001110010110100",
						 "100101101001110110001000",
						 "100101101001111001011100",
						 "100101101001111100110000",
						 "100101101010000000000100",
						 "100101101010000011011000",
						 "100101101010000110101100",
						 "100101101010001010000000",
						 "100101101010001101010100",
						 "100101101010010000101000",
						 "100101101010010011111100",
						 "100101101010010111010000",
						 "100101101001100101100100",
						 "100101101001101000111000",
						 "100101101001101100001100",
						 "100101101001101111100000",
						 "100101101001110010110100",
						 "100101101001110110001000",
						 "100101101001111001011100",
						 "100101101001111100110000",
						 "100101101010000000000100",
						 "100101101010000011011000",
						 "100101101010000110101100",
						 "100101101010001010000000",
						 "100101101010001101010100",
						 "100101101010010000101000",
						 "100101101010010011111100",
						 "100101101010010111010000",
						 "100101101001100101100100",
						 "100101101001101000110111",
						 "100101101001101100001010",
						 "100101101001101111011101",
						 "100101101001110010110000",
						 "100101101001110110000011",
						 "100101101001111001010110",
						 "100101101001111100101001",
						 "100101101001111111111100",
						 "100101101010000011001111",
						 "100101101010000110100010",
						 "100101101010001001110101",
						 "100101101010001101001000",
						 "100101101010010000011011",
						 "100101101010010011101110",
						 "100101101010010111000001",
						 "100101101100001000100010",
						 "100101101100001011110101",
						 "100101101100001111001000",
						 "100101101100010010011011",
						 "100101101100010101101110",
						 "100101101100011001000001",
						 "100101101100011100010100",
						 "100101101100011111100111",
						 "100101101100100010111010",
						 "100101101100100110001101",
						 "100101101100101001100000",
						 "100101101100101100110011",
						 "100101101100110000000110",
						 "100101101100110011011001",
						 "100101101100110110101100",
						 "100101101100111001111111",
						 "100101101100001000100010",
						 "100101101100001011110101",
						 "100101101100001111001000",
						 "100101101100010010011011",
						 "100101101100010101101110",
						 "100101101100011001000001",
						 "100101101100011100010100",
						 "100101101100011111100111",
						 "100101101100100010111010",
						 "100101101100100110001101",
						 "100101101100101001100000",
						 "100101101100101100110011",
						 "100101101100110000000110",
						 "100101101100110011011001",
						 "100101101100110110101100",
						 "100101101100111001111111",
						 "100101101100001000100010",
						 "100101101100001011110101",
						 "100101101100001111001000",
						 "100101101100010010011011",
						 "100101101100010101101110",
						 "100101101100011001000001",
						 "100101101100011100010100",
						 "100101101100011111100111",
						 "100101101100100010111010",
						 "100101101100100110001101",
						 "100101101100101001100000",
						 "100101101100101100110011",
						 "100101101100110000000110",
						 "100101101100110011011001",
						 "100101101100110110101100",
						 "100101101100111001111111",
						 "100101101110101011100000",
						 "100101101110101110110011",
						 "100101101110110010000110",
						 "100101101110110101011001",
						 "100101101110111000101100",
						 "100101101110111011111111",
						 "100101101110111111010010",
						 "100101101111000010100101",
						 "100101101111000101111000",
						 "100101101111001001001011",
						 "100101101111001100011110",
						 "100101101111001111110001",
						 "100101101111010011000100",
						 "100101101111010110010111",
						 "100101101111011001101010",
						 "100101101111011100111101",
						 "100101101110101011100000",
						 "100101101110101110110010",
						 "100101101110110010000100",
						 "100101101110110101010110",
						 "100101101110111000101000",
						 "100101101110111011111010",
						 "100101101110111111001100",
						 "100101101111000010011110",
						 "100101101111000101110000",
						 "100101101111001001000010",
						 "100101101111001100010100",
						 "100101101111001111100110",
						 "100101101111010010111000",
						 "100101101111010110001010",
						 "100101101111011001011100",
						 "100101101111011100101110",
						 "100101101110101011100000",
						 "100101101110101110110010",
						 "100101101110110010000100",
						 "100101101110110101010110",
						 "100101101110111000101000",
						 "100101101110111011111010",
						 "100101101110111111001100",
						 "100101101111000010011110",
						 "100101101111000101110000",
						 "100101101111001001000010",
						 "100101101111001100010100",
						 "100101101111001111100110",
						 "100101101111010010111000",
						 "100101101111010110001010",
						 "100101101111011001011100",
						 "100101101111011100101110",
						 "100101110001001110011110",
						 "100101110001010001110000",
						 "100101110001010101000010",
						 "100101110001011000010100",
						 "100101110001011011100110",
						 "100101110001011110111000",
						 "100101110001100010001010",
						 "100101110001100101011100",
						 "100101110001101000101110",
						 "100101110001101100000000",
						 "100101110001101111010010",
						 "100101110001110010100100",
						 "100101110001110101110110",
						 "100101110001111001001000",
						 "100101110001111100011010",
						 "100101110001111111101100",
						 "100101110001001110011110",
						 "100101110001010001110000",
						 "100101110001010101000010",
						 "100101110001011000010100",
						 "100101110001011011100110",
						 "100101110001011110111000",
						 "100101110001100010001010",
						 "100101110001100101011100",
						 "100101110001101000101110",
						 "100101110001101100000000",
						 "100101110001101111010010",
						 "100101110001110010100100",
						 "100101110001110101110110",
						 "100101110001111001001000",
						 "100101110001111100011010",
						 "100101110001111111101100",
						 "100101110001001110011110",
						 "100101110001010001101111",
						 "100101110001010101000000",
						 "100101110001011000010001",
						 "100101110001011011100010",
						 "100101110001011110110011",
						 "100101110001100010000100",
						 "100101110001100101010101",
						 "100101110001101000100110",
						 "100101110001101011110111",
						 "100101110001101111001000",
						 "100101110001110010011001",
						 "100101110001110101101010",
						 "100101110001111000111011",
						 "100101110001111100001100",
						 "100101110001111111011101",
						 "100101110011110001011100",
						 "100101110011110100101101",
						 "100101110011110111111110",
						 "100101110011111011001111",
						 "100101110011111110100000",
						 "100101110100000001110001",
						 "100101110100000101000010",
						 "100101110100001000010011",
						 "100101110100001011100100",
						 "100101110100001110110101",
						 "100101110100010010000110",
						 "100101110100010101010111",
						 "100101110100011000101000",
						 "100101110100011011111001",
						 "100101110100011111001010",
						 "100101110100100010011011",
						 "100101110011110001011100",
						 "100101110011110100101101",
						 "100101110011110111111110",
						 "100101110011111011001111",
						 "100101110011111110100000",
						 "100101110100000001110001",
						 "100101110100000101000010",
						 "100101110100001000010011",
						 "100101110100001011100100",
						 "100101110100001110110101",
						 "100101110100010010000110",
						 "100101110100010101010111",
						 "100101110100011000101000",
						 "100101110100011011111001",
						 "100101110100011111001010",
						 "100101110100100010011011",
						 "100101110011110001011100",
						 "100101110011110100101101",
						 "100101110011110111111110",
						 "100101110011111011001111",
						 "100101110011111110100000",
						 "100101110100000001110001",
						 "100101110100000101000010",
						 "100101110100001000010011",
						 "100101110100001011100100",
						 "100101110100001110110101",
						 "100101110100010010000110",
						 "100101110100010101010111",
						 "100101110100011000101000",
						 "100101110100011011111001",
						 "100101110100011111001010",
						 "100101110100100010011011",
						 "100101110110010100011010",
						 "100101110110010111101011",
						 "100101110110011010111100",
						 "100101110110011110001101",
						 "100101110110100001011110",
						 "100101110110100100101111",
						 "100101110110101000000000",
						 "100101110110101011010001",
						 "100101110110101110100010",
						 "100101110110110001110011",
						 "100101110110110101000100",
						 "100101110110111000010101",
						 "100101110110111011100110",
						 "100101110110111110110111",
						 "100101110111000010001000",
						 "100101110111000101011001",
						 "100101110110010100011010",
						 "100101110110010111101010",
						 "100101110110011010111010",
						 "100101110110011110001010",
						 "100101110110100001011010",
						 "100101110110100100101010",
						 "100101110110100111111010",
						 "100101110110101011001010",
						 "100101110110101110011010",
						 "100101110110110001101010",
						 "100101110110110100111010",
						 "100101110110111000001010",
						 "100101110110111011011010",
						 "100101110110111110101010",
						 "100101110111000001111010",
						 "100101110111000101001010",
						 "100101110110010100011010",
						 "100101110110010111101010",
						 "100101110110011010111010",
						 "100101110110011110001010",
						 "100101110110100001011010",
						 "100101110110100100101010",
						 "100101110110100111111010",
						 "100101110110101011001010",
						 "100101110110101110011010",
						 "100101110110110001101010",
						 "100101110110110100111010",
						 "100101110110111000001010",
						 "100101110110111011011010",
						 "100101110110111110101010",
						 "100101110111000001111010",
						 "100101110111000101001010",
						 "100101110110010100011010",
						 "100101110110010111101010",
						 "100101110110011010111010",
						 "100101110110011110001010",
						 "100101110110100001011010",
						 "100101110110100100101010",
						 "100101110110100111111010",
						 "100101110110101011001010",
						 "100101110110101110011010",
						 "100101110110110001101010",
						 "100101110110110100111010",
						 "100101110110111000001010",
						 "100101110110111011011010",
						 "100101110110111110101010",
						 "100101110111000001111010",
						 "100101110111000101001010",
						 "100101111000110111011000",
						 "100101111000111010101000",
						 "100101111000111101111000",
						 "100101111001000001001000",
						 "100101111001000100011000",
						 "100101111001000111101000",
						 "100101111001001010111000",
						 "100101111001001110001000",
						 "100101111001010001011000",
						 "100101111001010100101000",
						 "100101111001010111111000",
						 "100101111001011011001000",
						 "100101111001011110011000",
						 "100101111001100001101000",
						 "100101111001100100111000",
						 "100101111001101000001000",
						 "100101111000110111011000",
						 "100101111000111010100111",
						 "100101111000111101110110",
						 "100101111001000001000101",
						 "100101111001000100010100",
						 "100101111001000111100011",
						 "100101111001001010110010",
						 "100101111001001110000001",
						 "100101111001010001010000",
						 "100101111001010100011111",
						 "100101111001010111101110",
						 "100101111001011010111101",
						 "100101111001011110001100",
						 "100101111001100001011011",
						 "100101111001100100101010",
						 "100101111001100111111001",
						 "100101111000110111011000",
						 "100101111000111010100111",
						 "100101111000111101110110",
						 "100101111001000001000101",
						 "100101111001000100010100",
						 "100101111001000111100011",
						 "100101111001001010110010",
						 "100101111001001110000001",
						 "100101111001010001010000",
						 "100101111001010100011111",
						 "100101111001010111101110",
						 "100101111001011010111101",
						 "100101111001011110001100",
						 "100101111001100001011011",
						 "100101111001100100101010",
						 "100101111001100111111001",
						 "100101111011011010010110",
						 "100101111011011101100101",
						 "100101111011100000110100",
						 "100101111011100100000011",
						 "100101111011100111010010",
						 "100101111011101010100001",
						 "100101111011101101110000",
						 "100101111011110000111111",
						 "100101111011110100001110",
						 "100101111011110111011101",
						 "100101111011111010101100",
						 "100101111011111101111011",
						 "100101111100000001001010",
						 "100101111100000100011001",
						 "100101111100000111101000",
						 "100101111100001010110111",
						 "100101111011011010010110",
						 "100101111011011101100101",
						 "100101111011100000110100",
						 "100101111011100100000011",
						 "100101111011100111010010",
						 "100101111011101010100001",
						 "100101111011101101110000",
						 "100101111011110000111111",
						 "100101111011110100001110",
						 "100101111011110111011101",
						 "100101111011111010101100",
						 "100101111011111101111011",
						 "100101111100000001001010",
						 "100101111100000100011001",
						 "100101111100000111101000",
						 "100101111100001010110111",
						 "100101111011011010010110",
						 "100101111011011101100101",
						 "100101111011100000110100",
						 "100101111011100100000011",
						 "100101111011100111010010",
						 "100101111011101010100001",
						 "100101111011101101110000",
						 "100101111011110000111111",
						 "100101111011110100001110",
						 "100101111011110111011101",
						 "100101111011111010101100",
						 "100101111011111101111011",
						 "100101111100000001001010",
						 "100101111100000100011001",
						 "100101111100000111101000",
						 "100101111100001010110111",
						 "100101111101111101010100",
						 "100101111110000000100010",
						 "100101111110000011110000",
						 "100101111110000110111110",
						 "100101111110001010001100",
						 "100101111110001101011010",
						 "100101111110010000101000",
						 "100101111110010011110110",
						 "100101111110010111000100",
						 "100101111110011010010010",
						 "100101111110011101100000",
						 "100101111110100000101110",
						 "100101111110100011111100",
						 "100101111110100111001010",
						 "100101111110101010011000",
						 "100101111110101101100110",
						 "100101111101111101010100",
						 "100101111110000000100010",
						 "100101111110000011110000",
						 "100101111110000110111110",
						 "100101111110001010001100",
						 "100101111110001101011010",
						 "100101111110010000101000",
						 "100101111110010011110110",
						 "100101111110010111000100",
						 "100101111110011010010010",
						 "100101111110011101100000",
						 "100101111110100000101110",
						 "100101111110100011111100",
						 "100101111110100111001010",
						 "100101111110101010011000",
						 "100101111110101101100110",
						 "100101111101111101010100",
						 "100101111110000000100010",
						 "100101111110000011110000",
						 "100101111110000110111110",
						 "100101111110001010001100",
						 "100101111110001101011010",
						 "100101111110010000101000",
						 "100101111110010011110110",
						 "100101111110010111000100",
						 "100101111110011010010010",
						 "100101111110011101100000",
						 "100101111110100000101110",
						 "100101111110100011111100",
						 "100101111110100111001010",
						 "100101111110101010011000",
						 "100101111110101101100110",
						 "100110000000100000010010",
						 "100110000000100011100000",
						 "100110000000100110101110",
						 "100110000000101001111100",
						 "100110000000101101001010",
						 "100110000000110000011000",
						 "100110000000110011100110",
						 "100110000000110110110100",
						 "100110000000111010000010",
						 "100110000000111101010000",
						 "100110000001000000011110",
						 "100110000001000011101100",
						 "100110000001000110111010",
						 "100110000001001010001000",
						 "100110000001001101010110",
						 "100110000001010000100100",
						 "100110000000100000010010",
						 "100110000000100011011111",
						 "100110000000100110101100",
						 "100110000000101001111001",
						 "100110000000101101000110",
						 "100110000000110000010011",
						 "100110000000110011100000",
						 "100110000000110110101101",
						 "100110000000111001111010",
						 "100110000000111101000111",
						 "100110000001000000010100",
						 "100110000001000011100001",
						 "100110000001000110101110",
						 "100110000001001001111011",
						 "100110000001001101001000",
						 "100110000001010000010101",
						 "100110000000100000010010",
						 "100110000000100011011111",
						 "100110000000100110101100",
						 "100110000000101001111001",
						 "100110000000101101000110",
						 "100110000000110000010011",
						 "100110000000110011100000",
						 "100110000000110110101101",
						 "100110000000111001111010",
						 "100110000000111101000111",
						 "100110000001000000010100",
						 "100110000001000011100001",
						 "100110000001000110101110",
						 "100110000001001001111011",
						 "100110000001001101001000",
						 "100110000001010000010101",
						 "100110000011000011010000",
						 "100110000011000110011101",
						 "100110000011001001101010",
						 "100110000011001100110111",
						 "100110000011010000000100",
						 "100110000011010011010001",
						 "100110000011010110011110",
						 "100110000011011001101011",
						 "100110000011011100111000",
						 "100110000011100000000101",
						 "100110000011100011010010",
						 "100110000011100110011111",
						 "100110000011101001101100",
						 "100110000011101100111001",
						 "100110000011110000000110",
						 "100110000011110011010011",
						 "100110000011000011010000",
						 "100110000011000110011101",
						 "100110000011001001101010",
						 "100110000011001100110111",
						 "100110000011010000000100",
						 "100110000011010011010001",
						 "100110000011010110011110",
						 "100110000011011001101011",
						 "100110000011011100111000",
						 "100110000011100000000101",
						 "100110000011100011010010",
						 "100110000011100110011111",
						 "100110000011101001101100",
						 "100110000011101100111001",
						 "100110000011110000000110",
						 "100110000011110011010011",
						 "100110000011000011010000",
						 "100110000011000110011100",
						 "100110000011001001101000",
						 "100110000011001100110100",
						 "100110000011010000000000",
						 "100110000011010011001100",
						 "100110000011010110011000",
						 "100110000011011001100100",
						 "100110000011011100110000",
						 "100110000011011111111100",
						 "100110000011100011001000",
						 "100110000011100110010100",
						 "100110000011101001100000",
						 "100110000011101100101100",
						 "100110000011101111111000",
						 "100110000011110011000100",
						 "100110000101100110001110",
						 "100110000101101001011010",
						 "100110000101101100100110",
						 "100110000101101111110010",
						 "100110000101110010111110",
						 "100110000101110110001010",
						 "100110000101111001010110",
						 "100110000101111100100010",
						 "100110000101111111101110",
						 "100110000110000010111010",
						 "100110000110000110000110",
						 "100110000110001001010010",
						 "100110000110001100011110",
						 "100110000110001111101010",
						 "100110000110010010110110",
						 "100110000110010110000010",
						 "100110000101100110001110",
						 "100110000101101001011010",
						 "100110000101101100100110",
						 "100110000101101111110010",
						 "100110000101110010111110",
						 "100110000101110110001010",
						 "100110000101111001010110",
						 "100110000101111100100010",
						 "100110000101111111101110",
						 "100110000110000010111010",
						 "100110000110000110000110",
						 "100110000110001001010010",
						 "100110000110001100011110",
						 "100110000110001111101010",
						 "100110000110010010110110",
						 "100110000110010110000010",
						 "100110000101100110001110",
						 "100110000101101001011010",
						 "100110000101101100100110",
						 "100110000101101111110010",
						 "100110000101110010111110",
						 "100110000101110110001010",
						 "100110000101111001010110",
						 "100110000101111100100010",
						 "100110000101111111101110",
						 "100110000110000010111010",
						 "100110000110000110000110",
						 "100110000110001001010010",
						 "100110000110001100011110",
						 "100110000110001111101010",
						 "100110000110010010110110",
						 "100110000110010110000010",
						 "100110000101100110001110",
						 "100110000101101001011010",
						 "100110000101101100100110",
						 "100110000101101111110010",
						 "100110000101110010111110",
						 "100110000101110110001010",
						 "100110000101111001010110",
						 "100110000101111100100010",
						 "100110000101111111101110",
						 "100110000110000010111010",
						 "100110000110000110000110",
						 "100110000110001001010010",
						 "100110000110001100011110",
						 "100110000110001111101010",
						 "100110000110010010110110",
						 "100110000110010110000010",
						 "100110001000001001001100",
						 "100110001000001100010111",
						 "100110001000001111100010",
						 "100110001000010010101101",
						 "100110001000010101111000",
						 "100110001000011001000011",
						 "100110001000011100001110",
						 "100110001000011111011001",
						 "100110001000100010100100",
						 "100110001000100101101111",
						 "100110001000101000111010",
						 "100110001000101100000101",
						 "100110001000101111010000",
						 "100110001000110010011011",
						 "100110001000110101100110",
						 "100110001000111000110001",
						 "100110001000001001001100",
						 "100110001000001100010111",
						 "100110001000001111100010",
						 "100110001000010010101101",
						 "100110001000010101111000",
						 "100110001000011001000011",
						 "100110001000011100001110",
						 "100110001000011111011001",
						 "100110001000100010100100",
						 "100110001000100101101111",
						 "100110001000101000111010",
						 "100110001000101100000101",
						 "100110001000101111010000",
						 "100110001000110010011011",
						 "100110001000110101100110",
						 "100110001000111000110001",
						 "100110001000001001001100",
						 "100110001000001100010111",
						 "100110001000001111100010",
						 "100110001000010010101101",
						 "100110001000010101111000",
						 "100110001000011001000011",
						 "100110001000011100001110",
						 "100110001000011111011001",
						 "100110001000100010100100",
						 "100110001000100101101111",
						 "100110001000101000111010",
						 "100110001000101100000101",
						 "100110001000101111010000",
						 "100110001000110010011011",
						 "100110001000110101100110",
						 "100110001000111000110001",
						 "100110001010101100001010",
						 "100110001010101111010101",
						 "100110001010110010100000",
						 "100110001010110101101011",
						 "100110001010111000110110",
						 "100110001010111100000001",
						 "100110001010111111001100",
						 "100110001011000010010111",
						 "100110001011000101100010",
						 "100110001011001000101101",
						 "100110001011001011111000",
						 "100110001011001111000011",
						 "100110001011010010001110",
						 "100110001011010101011001",
						 "100110001011011000100100",
						 "100110001011011011101111",
						 "100110001010101100001010",
						 "100110001010101111010100",
						 "100110001010110010011110",
						 "100110001010110101101000",
						 "100110001010111000110010",
						 "100110001010111011111100",
						 "100110001010111111000110",
						 "100110001011000010010000",
						 "100110001011000101011010",
						 "100110001011001000100100",
						 "100110001011001011101110",
						 "100110001011001110111000",
						 "100110001011010010000010",
						 "100110001011010101001100",
						 "100110001011011000010110",
						 "100110001011011011100000",
						 "100110001010101100001010",
						 "100110001010101111010100",
						 "100110001010110010011110",
						 "100110001010110101101000",
						 "100110001010111000110010",
						 "100110001010111011111100",
						 "100110001010111111000110",
						 "100110001011000010010000",
						 "100110001011000101011010",
						 "100110001011001000100100",
						 "100110001011001011101110",
						 "100110001011001110111000",
						 "100110001011010010000010",
						 "100110001011010101001100",
						 "100110001011011000010110",
						 "100110001011011011100000",
						 "100110001101001111001000",
						 "100110001101010010010010",
						 "100110001101010101011100",
						 "100110001101011000100110",
						 "100110001101011011110000",
						 "100110001101011110111010",
						 "100110001101100010000100",
						 "100110001101100101001110",
						 "100110001101101000011000",
						 "100110001101101011100010",
						 "100110001101101110101100",
						 "100110001101110001110110",
						 "100110001101110101000000",
						 "100110001101111000001010",
						 "100110001101111011010100",
						 "100110001101111110011110",
						 "100110001101001111001000",
						 "100110001101010010010010",
						 "100110001101010101011100",
						 "100110001101011000100110",
						 "100110001101011011110000",
						 "100110001101011110111010",
						 "100110001101100010000100",
						 "100110001101100101001110",
						 "100110001101101000011000",
						 "100110001101101011100010",
						 "100110001101101110101100",
						 "100110001101110001110110",
						 "100110001101110101000000",
						 "100110001101111000001010",
						 "100110001101111011010100",
						 "100110001101111110011110",
						 "100110001101001111001000",
						 "100110001101010010010001",
						 "100110001101010101011010",
						 "100110001101011000100011",
						 "100110001101011011101100",
						 "100110001101011110110101",
						 "100110001101100001111110",
						 "100110001101100101000111",
						 "100110001101101000010000",
						 "100110001101101011011001",
						 "100110001101101110100010",
						 "100110001101110001101011",
						 "100110001101110100110100",
						 "100110001101110111111101",
						 "100110001101111011000110",
						 "100110001101111110001111",
						 "100110001111110010000110",
						 "100110001111110101001111",
						 "100110001111111000011000",
						 "100110001111111011100001",
						 "100110001111111110101010",
						 "100110010000000001110011",
						 "100110010000000100111100",
						 "100110010000001000000101",
						 "100110010000001011001110",
						 "100110010000001110010111",
						 "100110010000010001100000",
						 "100110010000010100101001",
						 "100110010000010111110010",
						 "100110010000011010111011",
						 "100110010000011110000100",
						 "100110010000100001001101",
						 "100110001111110010000110",
						 "100110001111110101001111",
						 "100110001111111000011000",
						 "100110001111111011100001",
						 "100110001111111110101010",
						 "100110010000000001110011",
						 "100110010000000100111100",
						 "100110010000001000000101",
						 "100110010000001011001110",
						 "100110010000001110010111",
						 "100110010000010001100000",
						 "100110010000010100101001",
						 "100110010000010111110010",
						 "100110010000011010111011",
						 "100110010000011110000100",
						 "100110010000100001001101",
						 "100110001111110010000110",
						 "100110001111110101001111",
						 "100110001111111000011000",
						 "100110001111111011100001",
						 "100110001111111110101010",
						 "100110010000000001110011",
						 "100110010000000100111100",
						 "100110010000001000000101",
						 "100110010000001011001110",
						 "100110010000001110010111",
						 "100110010000010001100000",
						 "100110010000010100101001",
						 "100110010000010111110010",
						 "100110010000011010111011",
						 "100110010000011110000100",
						 "100110010000100001001101",
						 "100110010010010101000100",
						 "100110010010011000001100",
						 "100110010010011011010100",
						 "100110010010011110011100",
						 "100110010010100001100100",
						 "100110010010100100101100",
						 "100110010010100111110100",
						 "100110010010101010111100",
						 "100110010010101110000100",
						 "100110010010110001001100",
						 "100110010010110100010100",
						 "100110010010110111011100",
						 "100110010010111010100100",
						 "100110010010111101101100",
						 "100110010011000000110100",
						 "100110010011000011111100",
						 "100110010010010101000100",
						 "100110010010011000001100",
						 "100110010010011011010100",
						 "100110010010011110011100",
						 "100110010010100001100100",
						 "100110010010100100101100",
						 "100110010010100111110100",
						 "100110010010101010111100",
						 "100110010010101110000100",
						 "100110010010110001001100",
						 "100110010010110100010100",
						 "100110010010110111011100",
						 "100110010010111010100100",
						 "100110010010111101101100",
						 "100110010011000000110100",
						 "100110010011000011111100",
						 "100110010010010101000100",
						 "100110010010011000001100",
						 "100110010010011011010100",
						 "100110010010011110011100",
						 "100110010010100001100100",
						 "100110010010100100101100",
						 "100110010010100111110100",
						 "100110010010101010111100",
						 "100110010010101110000100",
						 "100110010010110001001100",
						 "100110010010110100010100",
						 "100110010010110111011100",
						 "100110010010111010100100",
						 "100110010010111101101100",
						 "100110010011000000110100",
						 "100110010011000011111100",
						 "100110010010010101000100",
						 "100110010010011000001100",
						 "100110010010011011010100",
						 "100110010010011110011100",
						 "100110010010100001100100",
						 "100110010010100100101100",
						 "100110010010100111110100",
						 "100110010010101010111100",
						 "100110010010101110000100",
						 "100110010010110001001100",
						 "100110010010110100010100",
						 "100110010010110111011100",
						 "100110010010111010100100",
						 "100110010010111101101100",
						 "100110010011000000110100",
						 "100110010011000011111100",
						 "100110010100111000000010",
						 "100110010100111011001001",
						 "100110010100111110010000",
						 "100110010101000001010111",
						 "100110010101000100011110",
						 "100110010101000111100101",
						 "100110010101001010101100",
						 "100110010101001101110011",
						 "100110010101010000111010",
						 "100110010101010100000001",
						 "100110010101010111001000",
						 "100110010101011010001111",
						 "100110010101011101010110",
						 "100110010101100000011101",
						 "100110010101100011100100",
						 "100110010101100110101011",
						 "100110010100111000000010",
						 "100110010100111011001001",
						 "100110010100111110010000",
						 "100110010101000001010111",
						 "100110010101000100011110",
						 "100110010101000111100101",
						 "100110010101001010101100",
						 "100110010101001101110011",
						 "100110010101010000111010",
						 "100110010101010100000001",
						 "100110010101010111001000",
						 "100110010101011010001111",
						 "100110010101011101010110",
						 "100110010101100000011101",
						 "100110010101100011100100",
						 "100110010101100110101011",
						 "100110010100111000000010",
						 "100110010100111011001001",
						 "100110010100111110010000",
						 "100110010101000001010111",
						 "100110010101000100011110",
						 "100110010101000111100101",
						 "100110010101001010101100",
						 "100110010101001101110011",
						 "100110010101010000111010",
						 "100110010101010100000001",
						 "100110010101010111001000",
						 "100110010101011010001111",
						 "100110010101011101010110",
						 "100110010101100000011101",
						 "100110010101100011100100",
						 "100110010101100110101011",
						 "100110010111011011000000",
						 "100110010111011110000111",
						 "100110010111100001001110",
						 "100110010111100100010101",
						 "100110010111100111011100",
						 "100110010111101010100011",
						 "100110010111101101101010",
						 "100110010111110000110001",
						 "100110010111110011111000",
						 "100110010111110110111111",
						 "100110010111111010000110",
						 "100110010111111101001101",
						 "100110011000000000010100",
						 "100110011000000011011011",
						 "100110011000000110100010",
						 "100110011000001001101001",
						 "100110010111011011000000",
						 "100110010111011110000110",
						 "100110010111100001001100",
						 "100110010111100100010010",
						 "100110010111100111011000",
						 "100110010111101010011110",
						 "100110010111101101100100",
						 "100110010111110000101010",
						 "100110010111110011110000",
						 "100110010111110110110110",
						 "100110010111111001111100",
						 "100110010111111101000010",
						 "100110011000000000001000",
						 "100110011000000011001110",
						 "100110011000000110010100",
						 "100110011000001001011010",
						 "100110010111011011000000",
						 "100110010111011110000110",
						 "100110010111100001001100",
						 "100110010111100100010010",
						 "100110010111100111011000",
						 "100110010111101010011110",
						 "100110010111101101100100",
						 "100110010111110000101010",
						 "100110010111110011110000",
						 "100110010111110110110110",
						 "100110010111111001111100",
						 "100110010111111101000010",
						 "100110011000000000001000",
						 "100110011000000011001110",
						 "100110011000000110010100",
						 "100110011000001001011010",
						 "100110011001111101111110",
						 "100110011010000001000100",
						 "100110011010000100001010",
						 "100110011010000111010000",
						 "100110011010001010010110",
						 "100110011010001101011100",
						 "100110011010010000100010",
						 "100110011010010011101000",
						 "100110011010010110101110",
						 "100110011010011001110100",
						 "100110011010011100111010",
						 "100110011010100000000000",
						 "100110011010100011000110",
						 "100110011010100110001100",
						 "100110011010101001010010",
						 "100110011010101100011000",
						 "100110011001111101111110",
						 "100110011010000001000100",
						 "100110011010000100001010",
						 "100110011010000111010000",
						 "100110011010001010010110",
						 "100110011010001101011100",
						 "100110011010010000100010",
						 "100110011010010011101000",
						 "100110011010010110101110",
						 "100110011010011001110100",
						 "100110011010011100111010",
						 "100110011010100000000000",
						 "100110011010100011000110",
						 "100110011010100110001100",
						 "100110011010101001010010",
						 "100110011010101100011000",
						 "100110011001111101111110",
						 "100110011010000001000011",
						 "100110011010000100001000",
						 "100110011010000111001101",
						 "100110011010001010010010",
						 "100110011010001101010111",
						 "100110011010010000011100",
						 "100110011010010011100001",
						 "100110011010010110100110",
						 "100110011010011001101011",
						 "100110011010011100110000",
						 "100110011010011111110101",
						 "100110011010100010111010",
						 "100110011010100101111111",
						 "100110011010101001000100",
						 "100110011010101100001001",
						 "100110011001111101111110",
						 "100110011010000001000011",
						 "100110011010000100001000",
						 "100110011010000111001101",
						 "100110011010001010010010",
						 "100110011010001101010111",
						 "100110011010010000011100",
						 "100110011010010011100001",
						 "100110011010010110100110",
						 "100110011010011001101011",
						 "100110011010011100110000",
						 "100110011010011111110101",
						 "100110011010100010111010",
						 "100110011010100101111111",
						 "100110011010101001000100",
						 "100110011010101100001001",
						 "100110011100100000111100",
						 "100110011100100100000001",
						 "100110011100100111000110",
						 "100110011100101010001011",
						 "100110011100101101010000",
						 "100110011100110000010101",
						 "100110011100110011011010",
						 "100110011100110110011111",
						 "100110011100111001100100",
						 "100110011100111100101001",
						 "100110011100111111101110",
						 "100110011101000010110011",
						 "100110011101000101111000",
						 "100110011101001000111101",
						 "100110011101001100000010",
						 "100110011101001111000111",
						 "100110011100100000111100",
						 "100110011100100100000001",
						 "100110011100100111000110",
						 "100110011100101010001011",
						 "100110011100101101010000",
						 "100110011100110000010101",
						 "100110011100110011011010",
						 "100110011100110110011111",
						 "100110011100111001100100",
						 "100110011100111100101001",
						 "100110011100111111101110",
						 "100110011101000010110011",
						 "100110011101000101111000",
						 "100110011101001000111101",
						 "100110011101001100000010",
						 "100110011101001111000111",
						 "100110011100100000111100",
						 "100110011100100100000000",
						 "100110011100100111000100",
						 "100110011100101010001000",
						 "100110011100101101001100",
						 "100110011100110000010000",
						 "100110011100110011010100",
						 "100110011100110110011000",
						 "100110011100111001011100",
						 "100110011100111100100000",
						 "100110011100111111100100",
						 "100110011101000010101000",
						 "100110011101000101101100",
						 "100110011101001000110000",
						 "100110011101001011110100",
						 "100110011101001110111000",
						 "100110011111000011111010",
						 "100110011111000110111110",
						 "100110011111001010000010",
						 "100110011111001101000110",
						 "100110011111010000001010",
						 "100110011111010011001110",
						 "100110011111010110010010",
						 "100110011111011001010110",
						 "100110011111011100011010",
						 "100110011111011111011110",
						 "100110011111100010100010",
						 "100110011111100101100110",
						 "100110011111101000101010",
						 "100110011111101011101110",
						 "100110011111101110110010",
						 "100110011111110001110110",
						 "100110011111000011111010",
						 "100110011111000110111110",
						 "100110011111001010000010",
						 "100110011111001101000110",
						 "100110011111010000001010",
						 "100110011111010011001110",
						 "100110011111010110010010",
						 "100110011111011001010110",
						 "100110011111011100011010",
						 "100110011111011111011110",
						 "100110011111100010100010",
						 "100110011111100101100110",
						 "100110011111101000101010",
						 "100110011111101011101110",
						 "100110011111101110110010",
						 "100110011111110001110110",
						 "100110011111000011111010",
						 "100110011111000110111110",
						 "100110011111001010000010",
						 "100110011111001101000110",
						 "100110011111010000001010",
						 "100110011111010011001110",
						 "100110011111010110010010",
						 "100110011111011001010110",
						 "100110011111011100011010",
						 "100110011111011111011110",
						 "100110011111100010100010",
						 "100110011111100101100110",
						 "100110011111101000101010",
						 "100110011111101011101110",
						 "100110011111101110110010",
						 "100110011111110001110110",
						 "100110100001100110111000",
						 "100110100001101001111011",
						 "100110100001101100111110",
						 "100110100001110000000001",
						 "100110100001110011000100",
						 "100110100001110110000111",
						 "100110100001111001001010",
						 "100110100001111100001101",
						 "100110100001111111010000",
						 "100110100010000010010011",
						 "100110100010000101010110",
						 "100110100010001000011001",
						 "100110100010001011011100",
						 "100110100010001110011111",
						 "100110100010010001100010",
						 "100110100010010100100101",
						 "100110100001100110111000",
						 "100110100001101001111011",
						 "100110100001101100111110",
						 "100110100001110000000001",
						 "100110100001110011000100",
						 "100110100001110110000111",
						 "100110100001111001001010",
						 "100110100001111100001101",
						 "100110100001111111010000",
						 "100110100010000010010011",
						 "100110100010000101010110",
						 "100110100010001000011001",
						 "100110100010001011011100",
						 "100110100010001110011111",
						 "100110100010010001100010",
						 "100110100010010100100101",
						 "100110100001100110111000",
						 "100110100001101001111011",
						 "100110100001101100111110",
						 "100110100001110000000001",
						 "100110100001110011000100",
						 "100110100001110110000111",
						 "100110100001111001001010",
						 "100110100001111100001101",
						 "100110100001111111010000",
						 "100110100010000010010011",
						 "100110100010000101010110",
						 "100110100010001000011001",
						 "100110100010001011011100",
						 "100110100010001110011111",
						 "100110100010010001100010",
						 "100110100010010100100101",
						 "100110100001100110111000",
						 "100110100001101001111011",
						 "100110100001101100111110",
						 "100110100001110000000001",
						 "100110100001110011000100",
						 "100110100001110110000111",
						 "100110100001111001001010",
						 "100110100001111100001101",
						 "100110100001111111010000",
						 "100110100010000010010011",
						 "100110100010000101010110",
						 "100110100010001000011001",
						 "100110100010001011011100",
						 "100110100010001110011111",
						 "100110100010010001100010",
						 "100110100010010100100101",
						 "100110100100001001110110",
						 "100110100100001100111000",
						 "100110100100001111111010",
						 "100110100100010010111100",
						 "100110100100010101111110",
						 "100110100100011001000000",
						 "100110100100011100000010",
						 "100110100100011111000100",
						 "100110100100100010000110",
						 "100110100100100101001000",
						 "100110100100101000001010",
						 "100110100100101011001100",
						 "100110100100101110001110",
						 "100110100100110001010000",
						 "100110100100110100010010",
						 "100110100100110111010100",
						 "100110100100001001110110",
						 "100110100100001100111000",
						 "100110100100001111111010",
						 "100110100100010010111100",
						 "100110100100010101111110",
						 "100110100100011001000000",
						 "100110100100011100000010",
						 "100110100100011111000100",
						 "100110100100100010000110",
						 "100110100100100101001000",
						 "100110100100101000001010",
						 "100110100100101011001100",
						 "100110100100101110001110",
						 "100110100100110001010000",
						 "100110100100110100010010",
						 "100110100100110111010100",
						 "100110100100001001110110",
						 "100110100100001100111000",
						 "100110100100001111111010",
						 "100110100100010010111100",
						 "100110100100010101111110",
						 "100110100100011001000000",
						 "100110100100011100000010",
						 "100110100100011111000100",
						 "100110100100100010000110",
						 "100110100100100101001000",
						 "100110100100101000001010",
						 "100110100100101011001100",
						 "100110100100101110001110",
						 "100110100100110001010000",
						 "100110100100110100010010",
						 "100110100100110111010100",
						 "100110100110101100110100",
						 "100110100110101111110110",
						 "100110100110110010111000",
						 "100110100110110101111010",
						 "100110100110111000111100",
						 "100110100110111011111110",
						 "100110100110111111000000",
						 "100110100111000010000010",
						 "100110100111000101000100",
						 "100110100111001000000110",
						 "100110100111001011001000",
						 "100110100111001110001010",
						 "100110100111010001001100",
						 "100110100111010100001110",
						 "100110100111010111010000",
						 "100110100111011010010010",
						 "100110100110101100110100",
						 "100110100110101111110101",
						 "100110100110110010110110",
						 "100110100110110101110111",
						 "100110100110111000111000",
						 "100110100110111011111001",
						 "100110100110111110111010",
						 "100110100111000001111011",
						 "100110100111000100111100",
						 "100110100111000111111101",
						 "100110100111001010111110",
						 "100110100111001101111111",
						 "100110100111010001000000",
						 "100110100111010100000001",
						 "100110100111010111000010",
						 "100110100111011010000011",
						 "100110100110101100110100",
						 "100110100110101111110101",
						 "100110100110110010110110",
						 "100110100110110101110111",
						 "100110100110111000111000",
						 "100110100110111011111001",
						 "100110100110111110111010",
						 "100110100111000001111011",
						 "100110100111000100111100",
						 "100110100111000111111101",
						 "100110100111001010111110",
						 "100110100111001101111111",
						 "100110100111010001000000",
						 "100110100111010100000001",
						 "100110100111010111000010",
						 "100110100111011010000011",
						 "100110101001001111110010",
						 "100110101001010010110011",
						 "100110101001010101110100",
						 "100110101001011000110101",
						 "100110101001011011110110",
						 "100110101001011110110111",
						 "100110101001100001111000",
						 "100110101001100100111001",
						 "100110101001100111111010",
						 "100110101001101010111011",
						 "100110101001101101111100",
						 "100110101001110000111101",
						 "100110101001110011111110",
						 "100110101001110110111111",
						 "100110101001111010000000",
						 "100110101001111101000001",
						 "100110101001001111110010",
						 "100110101001010010110011",
						 "100110101001010101110100",
						 "100110101001011000110101",
						 "100110101001011011110110",
						 "100110101001011110110111",
						 "100110101001100001111000",
						 "100110101001100100111001",
						 "100110101001100111111010",
						 "100110101001101010111011",
						 "100110101001101101111100",
						 "100110101001110000111101",
						 "100110101001110011111110",
						 "100110101001110110111111",
						 "100110101001111010000000",
						 "100110101001111101000001",
						 "100110101001001111110010",
						 "100110101001010010110010",
						 "100110101001010101110010",
						 "100110101001011000110010",
						 "100110101001011011110010",
						 "100110101001011110110010",
						 "100110101001100001110010",
						 "100110101001100100110010",
						 "100110101001100111110010",
						 "100110101001101010110010",
						 "100110101001101101110010",
						 "100110101001110000110010",
						 "100110101001110011110010",
						 "100110101001110110110010",
						 "100110101001111001110010",
						 "100110101001111100110010",
						 "100110101001001111110010",
						 "100110101001010010110010",
						 "100110101001010101110010",
						 "100110101001011000110010",
						 "100110101001011011110010",
						 "100110101001011110110010",
						 "100110101001100001110010",
						 "100110101001100100110010",
						 "100110101001100111110010",
						 "100110101001101010110010",
						 "100110101001101101110010",
						 "100110101001110000110010",
						 "100110101001110011110010",
						 "100110101001110110110010",
						 "100110101001111001110010",
						 "100110101001111100110010",
						 "100110101011110010110000",
						 "100110101011110101110000",
						 "100110101011111000110000",
						 "100110101011111011110000",
						 "100110101011111110110000",
						 "100110101100000001110000",
						 "100110101100000100110000",
						 "100110101100000111110000",
						 "100110101100001010110000",
						 "100110101100001101110000",
						 "100110101100010000110000",
						 "100110101100010011110000",
						 "100110101100010110110000",
						 "100110101100011001110000",
						 "100110101100011100110000",
						 "100110101100011111110000",
						 "100110101011110010110000",
						 "100110101011110101110000",
						 "100110101011111000110000",
						 "100110101011111011110000",
						 "100110101011111110110000",
						 "100110101100000001110000",
						 "100110101100000100110000",
						 "100110101100000111110000",
						 "100110101100001010110000",
						 "100110101100001101110000",
						 "100110101100010000110000",
						 "100110101100010011110000",
						 "100110101100010110110000",
						 "100110101100011001110000",
						 "100110101100011100110000",
						 "100110101100011111110000",
						 "100110101011110010110000",
						 "100110101011110101101111",
						 "100110101011111000101110",
						 "100110101011111011101101",
						 "100110101011111110101100",
						 "100110101100000001101011",
						 "100110101100000100101010",
						 "100110101100000111101001",
						 "100110101100001010101000",
						 "100110101100001101100111",
						 "100110101100010000100110",
						 "100110101100010011100101",
						 "100110101100010110100100",
						 "100110101100011001100011",
						 "100110101100011100100010",
						 "100110101100011111100001",
						 "100110101110010101101110",
						 "100110101110011000101101",
						 "100110101110011011101100",
						 "100110101110011110101011",
						 "100110101110100001101010",
						 "100110101110100100101001",
						 "100110101110100111101000",
						 "100110101110101010100111",
						 "100110101110101101100110",
						 "100110101110110000100101",
						 "100110101110110011100100",
						 "100110101110110110100011",
						 "100110101110111001100010",
						 "100110101110111100100001",
						 "100110101110111111100000",
						 "100110101111000010011111",
						 "100110101110010101101110",
						 "100110101110011000101101",
						 "100110101110011011101100",
						 "100110101110011110101011",
						 "100110101110100001101010",
						 "100110101110100100101001",
						 "100110101110100111101000",
						 "100110101110101010100111",
						 "100110101110101101100110",
						 "100110101110110000100101",
						 "100110101110110011100100",
						 "100110101110110110100011",
						 "100110101110111001100010",
						 "100110101110111100100001",
						 "100110101110111111100000",
						 "100110101111000010011111",
						 "100110101110010101101110",
						 "100110101110011000101101",
						 "100110101110011011101100",
						 "100110101110011110101011",
						 "100110101110100001101010",
						 "100110101110100100101001",
						 "100110101110100111101000",
						 "100110101110101010100111",
						 "100110101110101101100110",
						 "100110101110110000100101",
						 "100110101110110011100100",
						 "100110101110110110100011",
						 "100110101110111001100010",
						 "100110101110111100100001",
						 "100110101110111111100000",
						 "100110101111000010011111",
						 "100110110000111000101100",
						 "100110110000111011101010",
						 "100110110000111110101000",
						 "100110110001000001100110",
						 "100110110001000100100100",
						 "100110110001000111100010",
						 "100110110001001010100000",
						 "100110110001001101011110",
						 "100110110001010000011100",
						 "100110110001010011011010",
						 "100110110001010110011000",
						 "100110110001011001010110",
						 "100110110001011100010100",
						 "100110110001011111010010",
						 "100110110001100010010000",
						 "100110110001100101001110",
						 "100110110000111000101100",
						 "100110110000111011101010",
						 "100110110000111110101000",
						 "100110110001000001100110",
						 "100110110001000100100100",
						 "100110110001000111100010",
						 "100110110001001010100000",
						 "100110110001001101011110",
						 "100110110001010000011100",
						 "100110110001010011011010",
						 "100110110001010110011000",
						 "100110110001011001010110",
						 "100110110001011100010100",
						 "100110110001011111010010",
						 "100110110001100010010000",
						 "100110110001100101001110",
						 "100110110000111000101100",
						 "100110110000111011101010",
						 "100110110000111110101000",
						 "100110110001000001100110",
						 "100110110001000100100100",
						 "100110110001000111100010",
						 "100110110001001010100000",
						 "100110110001001101011110",
						 "100110110001010000011100",
						 "100110110001010011011010",
						 "100110110001010110011000",
						 "100110110001011001010110",
						 "100110110001011100010100",
						 "100110110001011111010010",
						 "100110110001100010010000",
						 "100110110001100101001110",
						 "100110110000111000101100",
						 "100110110000111011101010",
						 "100110110000111110101000",
						 "100110110001000001100110",
						 "100110110001000100100100",
						 "100110110001000111100010",
						 "100110110001001010100000",
						 "100110110001001101011110",
						 "100110110001010000011100",
						 "100110110001010011011010",
						 "100110110001010110011000",
						 "100110110001011001010110",
						 "100110110001011100010100",
						 "100110110001011111010010",
						 "100110110001100010010000",
						 "100110110001100101001110",
						 "100110110011011011101010",
						 "100110110011011110100111",
						 "100110110011100001100100",
						 "100110110011100100100001",
						 "100110110011100111011110",
						 "100110110011101010011011",
						 "100110110011101101011000",
						 "100110110011110000010101",
						 "100110110011110011010010",
						 "100110110011110110001111",
						 "100110110011111001001100",
						 "100110110011111100001001",
						 "100110110011111111000110",
						 "100110110100000010000011",
						 "100110110100000101000000",
						 "100110110100000111111101",
						 "100110110011011011101010",
						 "100110110011011110100111",
						 "100110110011100001100100",
						 "100110110011100100100001",
						 "100110110011100111011110",
						 "100110110011101010011011",
						 "100110110011101101011000",
						 "100110110011110000010101",
						 "100110110011110011010010",
						 "100110110011110110001111",
						 "100110110011111001001100",
						 "100110110011111100001001",
						 "100110110011111111000110",
						 "100110110100000010000011",
						 "100110110100000101000000",
						 "100110110100000111111101",
						 "100110110011011011101010",
						 "100110110011011110100111",
						 "100110110011100001100100",
						 "100110110011100100100001",
						 "100110110011100111011110",
						 "100110110011101010011011",
						 "100110110011101101011000",
						 "100110110011110000010101",
						 "100110110011110011010010",
						 "100110110011110110001111",
						 "100110110011111001001100",
						 "100110110011111100001001",
						 "100110110011111111000110",
						 "100110110100000010000011",
						 "100110110100000101000000",
						 "100110110100000111111101",
						 "100110110101111110101000",
						 "100110110110000001100101",
						 "100110110110000100100010",
						 "100110110110000111011111",
						 "100110110110001010011100",
						 "100110110110001101011001",
						 "100110110110010000010110",
						 "100110110110010011010011",
						 "100110110110010110010000",
						 "100110110110011001001101",
						 "100110110110011100001010",
						 "100110110110011111000111",
						 "100110110110100010000100",
						 "100110110110100101000001",
						 "100110110110100111111110",
						 "100110110110101010111011",
						 "100110110101111110101000",
						 "100110110110000001100100",
						 "100110110110000100100000",
						 "100110110110000111011100",
						 "100110110110001010011000",
						 "100110110110001101010100",
						 "100110110110010000010000",
						 "100110110110010011001100",
						 "100110110110010110001000",
						 "100110110110011001000100",
						 "100110110110011100000000",
						 "100110110110011110111100",
						 "100110110110100001111000",
						 "100110110110100100110100",
						 "100110110110100111110000",
						 "100110110110101010101100",
						 "100110110101111110101000",
						 "100110110110000001100100",
						 "100110110110000100100000",
						 "100110110110000111011100",
						 "100110110110001010011000",
						 "100110110110001101010100",
						 "100110110110010000010000",
						 "100110110110010011001100",
						 "100110110110010110001000",
						 "100110110110011001000100",
						 "100110110110011100000000",
						 "100110110110011110111100",
						 "100110110110100001111000",
						 "100110110110100100110100",
						 "100110110110100111110000",
						 "100110110110101010101100",
						 "100110110101111110101000",
						 "100110110110000001100100",
						 "100110110110000100100000",
						 "100110110110000111011100",
						 "100110110110001010011000",
						 "100110110110001101010100",
						 "100110110110010000010000",
						 "100110110110010011001100",
						 "100110110110010110001000",
						 "100110110110011001000100",
						 "100110110110011100000000",
						 "100110110110011110111100",
						 "100110110110100001111000",
						 "100110110110100100110100",
						 "100110110110100111110000",
						 "100110110110101010101100",
						 "100110111000100001100110",
						 "100110111000100100100001",
						 "100110111000100111011100",
						 "100110111000101010010111",
						 "100110111000101101010010",
						 "100110111000110000001101",
						 "100110111000110011001000",
						 "100110111000110110000011",
						 "100110111000111000111110",
						 "100110111000111011111001",
						 "100110111000111110110100",
						 "100110111001000001101111",
						 "100110111001000100101010",
						 "100110111001000111100101",
						 "100110111001001010100000",
						 "100110111001001101011011",
						 "100110111000100001100110",
						 "100110111000100100100001",
						 "100110111000100111011100",
						 "100110111000101010010111",
						 "100110111000101101010010",
						 "100110111000110000001101",
						 "100110111000110011001000",
						 "100110111000110110000011",
						 "100110111000111000111110",
						 "100110111000111011111001",
						 "100110111000111110110100",
						 "100110111001000001101111",
						 "100110111001000100101010",
						 "100110111001000111100101",
						 "100110111001001010100000",
						 "100110111001001101011011",
						 "100110111000100001100110",
						 "100110111000100100100001",
						 "100110111000100111011100",
						 "100110111000101010010111",
						 "100110111000101101010010",
						 "100110111000110000001101",
						 "100110111000110011001000",
						 "100110111000110110000011",
						 "100110111000111000111110",
						 "100110111000111011111001",
						 "100110111000111110110100",
						 "100110111001000001101111",
						 "100110111001000100101010",
						 "100110111001000111100101",
						 "100110111001001010100000",
						 "100110111001001101011011",
						 "100110111011000100100100",
						 "100110111011000111011111",
						 "100110111011001010011010",
						 "100110111011001101010101",
						 "100110111011010000010000",
						 "100110111011010011001011",
						 "100110111011010110000110",
						 "100110111011011001000001",
						 "100110111011011011111100",
						 "100110111011011110110111",
						 "100110111011100001110010",
						 "100110111011100100101101",
						 "100110111011100111101000",
						 "100110111011101010100011",
						 "100110111011101101011110",
						 "100110111011110000011001",
						 "100110111011000100100100",
						 "100110111011000111011110",
						 "100110111011001010011000",
						 "100110111011001101010010",
						 "100110111011010000001100",
						 "100110111011010011000110",
						 "100110111011010110000000",
						 "100110111011011000111010",
						 "100110111011011011110100",
						 "100110111011011110101110",
						 "100110111011100001101000",
						 "100110111011100100100010",
						 "100110111011100111011100",
						 "100110111011101010010110",
						 "100110111011101101010000",
						 "100110111011110000001010",
						 "100110111011000100100100",
						 "100110111011000111011110",
						 "100110111011001010011000",
						 "100110111011001101010010",
						 "100110111011010000001100",
						 "100110111011010011000110",
						 "100110111011010110000000",
						 "100110111011011000111010",
						 "100110111011011011110100",
						 "100110111011011110101110",
						 "100110111011100001101000",
						 "100110111011100100100010",
						 "100110111011100111011100",
						 "100110111011101010010110",
						 "100110111011101101010000",
						 "100110111011110000001010",
						 "100110111011000100100100",
						 "100110111011000111011110",
						 "100110111011001010011000",
						 "100110111011001101010010",
						 "100110111011010000001100",
						 "100110111011010011000110",
						 "100110111011010110000000",
						 "100110111011011000111010",
						 "100110111011011011110100",
						 "100110111011011110101110",
						 "100110111011100001101000",
						 "100110111011100100100010",
						 "100110111011100111011100",
						 "100110111011101010010110",
						 "100110111011101101010000",
						 "100110111011110000001010",
						 "100110111101100111100010",
						 "100110111101101010011100",
						 "100110111101101101010110",
						 "100110111101110000010000",
						 "100110111101110011001010",
						 "100110111101110110000100",
						 "100110111101111000111110",
						 "100110111101111011111000",
						 "100110111101111110110010",
						 "100110111110000001101100",
						 "100110111110000100100110",
						 "100110111110000111100000",
						 "100110111110001010011010",
						 "100110111110001101010100",
						 "100110111110010000001110",
						 "100110111110010011001000",
						 "100110111101100111100010",
						 "100110111101101010011011",
						 "100110111101101101010100",
						 "100110111101110000001101",
						 "100110111101110011000110",
						 "100110111101110101111111",
						 "100110111101111000111000",
						 "100110111101111011110001",
						 "100110111101111110101010",
						 "100110111110000001100011",
						 "100110111110000100011100",
						 "100110111110000111010101",
						 "100110111110001010001110",
						 "100110111110001101000111",
						 "100110111110010000000000",
						 "100110111110010010111001",
						 "100110111101100111100010",
						 "100110111101101010011011",
						 "100110111101101101010100",
						 "100110111101110000001101",
						 "100110111101110011000110",
						 "100110111101110101111111",
						 "100110111101111000111000",
						 "100110111101111011110001",
						 "100110111101111110101010",
						 "100110111110000001100011",
						 "100110111110000100011100",
						 "100110111110000111010101",
						 "100110111110001010001110",
						 "100110111110001101000111",
						 "100110111110010000000000",
						 "100110111110010010111001",
						 "100111000000001010100000",
						 "100111000000001101011001",
						 "100111000000010000010010",
						 "100111000000010011001011",
						 "100111000000010110000100",
						 "100111000000011000111101",
						 "100111000000011011110110",
						 "100111000000011110101111",
						 "100111000000100001101000",
						 "100111000000100100100001",
						 "100111000000100111011010",
						 "100111000000101010010011",
						 "100111000000101101001100",
						 "100111000000110000000101",
						 "100111000000110010111110",
						 "100111000000110101110111",
						 "100111000000001010100000",
						 "100111000000001101011001",
						 "100111000000010000010010",
						 "100111000000010011001011",
						 "100111000000010110000100",
						 "100111000000011000111101",
						 "100111000000011011110110",
						 "100111000000011110101111",
						 "100111000000100001101000",
						 "100111000000100100100001",
						 "100111000000100111011010",
						 "100111000000101010010011",
						 "100111000000101101001100",
						 "100111000000110000000101",
						 "100111000000110010111110",
						 "100111000000110101110111",
						 "100111000000001010100000",
						 "100111000000001101011000",
						 "100111000000010000010000",
						 "100111000000010011001000",
						 "100111000000010110000000",
						 "100111000000011000111000",
						 "100111000000011011110000",
						 "100111000000011110101000",
						 "100111000000100001100000",
						 "100111000000100100011000",
						 "100111000000100111010000",
						 "100111000000101010001000",
						 "100111000000101101000000",
						 "100111000000101111111000",
						 "100111000000110010110000",
						 "100111000000110101101000",
						 "100111000000001010100000",
						 "100111000000001101011000",
						 "100111000000010000010000",
						 "100111000000010011001000",
						 "100111000000010110000000",
						 "100111000000011000111000",
						 "100111000000011011110000",
						 "100111000000011110101000",
						 "100111000000100001100000",
						 "100111000000100100011000",
						 "100111000000100111010000",
						 "100111000000101010001000",
						 "100111000000101101000000",
						 "100111000000101111111000",
						 "100111000000110010110000",
						 "100111000000110101101000",
						 "100111000010101101011110",
						 "100111000010110000010110",
						 "100111000010110011001110",
						 "100111000010110110000110",
						 "100111000010111000111110",
						 "100111000010111011110110",
						 "100111000010111110101110",
						 "100111000011000001100110",
						 "100111000011000100011110",
						 "100111000011000111010110",
						 "100111000011001010001110",
						 "100111000011001101000110",
						 "100111000011001111111110",
						 "100111000011010010110110",
						 "100111000011010101101110",
						 "100111000011011000100110",
						 "100111000010101101011110",
						 "100111000010110000010101",
						 "100111000010110011001100",
						 "100111000010110110000011",
						 "100111000010111000111010",
						 "100111000010111011110001",
						 "100111000010111110101000",
						 "100111000011000001011111",
						 "100111000011000100010110",
						 "100111000011000111001101",
						 "100111000011001010000100",
						 "100111000011001100111011",
						 "100111000011001111110010",
						 "100111000011010010101001",
						 "100111000011010101100000",
						 "100111000011011000010111",
						 "100111000010101101011110",
						 "100111000010110000010101",
						 "100111000010110011001100",
						 "100111000010110110000011",
						 "100111000010111000111010",
						 "100111000010111011110001",
						 "100111000010111110101000",
						 "100111000011000001011111",
						 "100111000011000100010110",
						 "100111000011000111001101",
						 "100111000011001010000100",
						 "100111000011001100111011",
						 "100111000011001111110010",
						 "100111000011010010101001",
						 "100111000011010101100000",
						 "100111000011011000010111",
						 "100111000101010000011100",
						 "100111000101010011010011",
						 "100111000101010110001010",
						 "100111000101011001000001",
						 "100111000101011011111000",
						 "100111000101011110101111",
						 "100111000101100001100110",
						 "100111000101100100011101",
						 "100111000101100111010100",
						 "100111000101101010001011",
						 "100111000101101101000010",
						 "100111000101101111111001",
						 "100111000101110010110000",
						 "100111000101110101100111",
						 "100111000101111000011110",
						 "100111000101111011010101",
						 "100111000101010000011100",
						 "100111000101010011010011",
						 "100111000101010110001010",
						 "100111000101011001000001",
						 "100111000101011011111000",
						 "100111000101011110101111",
						 "100111000101100001100110",
						 "100111000101100100011101",
						 "100111000101100111010100",
						 "100111000101101010001011",
						 "100111000101101101000010",
						 "100111000101101111111001",
						 "100111000101110010110000",
						 "100111000101110101100111",
						 "100111000101111000011110",
						 "100111000101111011010101",
						 "100111000101010000011100",
						 "100111000101010011010010",
						 "100111000101010110001000",
						 "100111000101011000111110",
						 "100111000101011011110100",
						 "100111000101011110101010",
						 "100111000101100001100000",
						 "100111000101100100010110",
						 "100111000101100111001100",
						 "100111000101101010000010",
						 "100111000101101100111000",
						 "100111000101101111101110",
						 "100111000101110010100100",
						 "100111000101110101011010",
						 "100111000101111000010000",
						 "100111000101111011000110",
						 "100111000101010000011100",
						 "100111000101010011010010",
						 "100111000101010110001000",
						 "100111000101011000111110",
						 "100111000101011011110100",
						 "100111000101011110101010",
						 "100111000101100001100000",
						 "100111000101100100010110",
						 "100111000101100111001100",
						 "100111000101101010000010",
						 "100111000101101100111000",
						 "100111000101101111101110",
						 "100111000101110010100100",
						 "100111000101110101011010",
						 "100111000101111000010000",
						 "100111000101111011000110",
						 "100111000111110011011010",
						 "100111000111110110010000",
						 "100111000111111001000110",
						 "100111000111111011111100",
						 "100111000111111110110010",
						 "100111001000000001101000",
						 "100111001000000100011110",
						 "100111001000000111010100",
						 "100111001000001010001010",
						 "100111001000001101000000",
						 "100111001000001111110110",
						 "100111001000010010101100",
						 "100111001000010101100010",
						 "100111001000011000011000",
						 "100111001000011011001110",
						 "100111001000011110000100",
						 "100111000111110011011010",
						 "100111000111110110010000",
						 "100111000111111001000110",
						 "100111000111111011111100",
						 "100111000111111110110010",
						 "100111001000000001101000",
						 "100111001000000100011110",
						 "100111001000000111010100",
						 "100111001000001010001010",
						 "100111001000001101000000",
						 "100111001000001111110110",
						 "100111001000010010101100",
						 "100111001000010101100010",
						 "100111001000011000011000",
						 "100111001000011011001110",
						 "100111001000011110000100",
						 "100111000111110011011010",
						 "100111000111110110001111",
						 "100111000111111001000100",
						 "100111000111111011111001",
						 "100111000111111110101110",
						 "100111001000000001100011",
						 "100111001000000100011000",
						 "100111001000000111001101",
						 "100111001000001010000010",
						 "100111001000001100110111",
						 "100111001000001111101100",
						 "100111001000010010100001",
						 "100111001000010101010110",
						 "100111001000011000001011",
						 "100111001000011011000000",
						 "100111001000011101110101",
						 "100111000111110011011010",
						 "100111000111110110001111",
						 "100111000111111001000100",
						 "100111000111111011111001",
						 "100111000111111110101110",
						 "100111001000000001100011",
						 "100111001000000100011000",
						 "100111001000000111001101",
						 "100111001000001010000010",
						 "100111001000001100110111",
						 "100111001000001111101100",
						 "100111001000010010100001",
						 "100111001000010101010110",
						 "100111001000011000001011",
						 "100111001000011011000000",
						 "100111001000011101110101",
						 "100111001010010110011000",
						 "100111001010011001001101",
						 "100111001010011100000010",
						 "100111001010011110110111",
						 "100111001010100001101100",
						 "100111001010100100100001",
						 "100111001010100111010110",
						 "100111001010101010001011",
						 "100111001010101101000000",
						 "100111001010101111110101",
						 "100111001010110010101010",
						 "100111001010110101011111",
						 "100111001010111000010100",
						 "100111001010111011001001",
						 "100111001010111101111110",
						 "100111001011000000110011",
						 "100111001010010110011000",
						 "100111001010011001001100",
						 "100111001010011100000000",
						 "100111001010011110110100",
						 "100111001010100001101000",
						 "100111001010100100011100",
						 "100111001010100111010000",
						 "100111001010101010000100",
						 "100111001010101100111000",
						 "100111001010101111101100",
						 "100111001010110010100000",
						 "100111001010110101010100",
						 "100111001010111000001000",
						 "100111001010111010111100",
						 "100111001010111101110000",
						 "100111001011000000100100",
						 "100111001010010110011000",
						 "100111001010011001001100",
						 "100111001010011100000000",
						 "100111001010011110110100",
						 "100111001010100001101000",
						 "100111001010100100011100",
						 "100111001010100111010000",
						 "100111001010101010000100",
						 "100111001010101100111000",
						 "100111001010101111101100",
						 "100111001010110010100000",
						 "100111001010110101010100",
						 "100111001010111000001000",
						 "100111001010111010111100",
						 "100111001010111101110000",
						 "100111001011000000100100",
						 "100111001100111001010110",
						 "100111001100111100001010",
						 "100111001100111110111110",
						 "100111001101000001110010",
						 "100111001101000100100110",
						 "100111001101000111011010",
						 "100111001101001010001110",
						 "100111001101001101000010",
						 "100111001101001111110110",
						 "100111001101010010101010",
						 "100111001101010101011110",
						 "100111001101011000010010",
						 "100111001101011011000110",
						 "100111001101011101111010",
						 "100111001101100000101110",
						 "100111001101100011100010",
						 "100111001100111001010110",
						 "100111001100111100001010",
						 "100111001100111110111110",
						 "100111001101000001110010",
						 "100111001101000100100110",
						 "100111001101000111011010",
						 "100111001101001010001110",
						 "100111001101001101000010",
						 "100111001101001111110110",
						 "100111001101010010101010",
						 "100111001101010101011110",
						 "100111001101011000010010",
						 "100111001101011011000110",
						 "100111001101011101111010",
						 "100111001101100000101110",
						 "100111001101100011100010",
						 "100111001100111001010110",
						 "100111001100111100001001",
						 "100111001100111110111100",
						 "100111001101000001101111",
						 "100111001101000100100010",
						 "100111001101000111010101",
						 "100111001101001010001000",
						 "100111001101001100111011",
						 "100111001101001111101110",
						 "100111001101010010100001",
						 "100111001101010101010100",
						 "100111001101011000000111",
						 "100111001101011010111010",
						 "100111001101011101101101",
						 "100111001101100000100000",
						 "100111001101100011010011",
						 "100111001100111001010110",
						 "100111001100111100001001",
						 "100111001100111110111100",
						 "100111001101000001101111",
						 "100111001101000100100010",
						 "100111001101000111010101",
						 "100111001101001010001000",
						 "100111001101001100111011",
						 "100111001101001111101110",
						 "100111001101010010100001",
						 "100111001101010101010100",
						 "100111001101011000000111",
						 "100111001101011010111010",
						 "100111001101011101101101",
						 "100111001101100000100000",
						 "100111001101100011010011",
						 "100111001111011100010100",
						 "100111001111011111000111",
						 "100111001111100001111010",
						 "100111001111100100101101",
						 "100111001111100111100000",
						 "100111001111101010010011",
						 "100111001111101101000110",
						 "100111001111101111111001",
						 "100111001111110010101100",
						 "100111001111110101011111",
						 "100111001111111000010010",
						 "100111001111111011000101",
						 "100111001111111101111000",
						 "100111010000000000101011",
						 "100111010000000011011110",
						 "100111010000000110010001",
						 "100111001111011100010100",
						 "100111001111011111000111",
						 "100111001111100001111010",
						 "100111001111100100101101",
						 "100111001111100111100000",
						 "100111001111101010010011",
						 "100111001111101101000110",
						 "100111001111101111111001",
						 "100111001111110010101100",
						 "100111001111110101011111",
						 "100111001111111000010010",
						 "100111001111111011000101",
						 "100111001111111101111000",
						 "100111010000000000101011",
						 "100111010000000011011110",
						 "100111010000000110010001",
						 "100111001111011100010100",
						 "100111001111011111000110",
						 "100111001111100001111000",
						 "100111001111100100101010",
						 "100111001111100111011100",
						 "100111001111101010001110",
						 "100111001111101101000000",
						 "100111001111101111110010",
						 "100111001111110010100100",
						 "100111001111110101010110",
						 "100111001111111000001000",
						 "100111001111111010111010",
						 "100111001111111101101100",
						 "100111010000000000011110",
						 "100111010000000011010000",
						 "100111010000000110000010",
						 "100111010001111111010010",
						 "100111010010000010000100",
						 "100111010010000100110110",
						 "100111010010000111101000",
						 "100111010010001010011010",
						 "100111010010001101001100",
						 "100111010010001111111110",
						 "100111010010010010110000",
						 "100111010010010101100010",
						 "100111010010011000010100",
						 "100111010010011011000110",
						 "100111010010011101111000",
						 "100111010010100000101010",
						 "100111010010100011011100",
						 "100111010010100110001110",
						 "100111010010101001000000",
						 "100111010001111111010010",
						 "100111010010000010000100",
						 "100111010010000100110110",
						 "100111010010000111101000",
						 "100111010010001010011010",
						 "100111010010001101001100",
						 "100111010010001111111110",
						 "100111010010010010110000",
						 "100111010010010101100010",
						 "100111010010011000010100",
						 "100111010010011011000110",
						 "100111010010011101111000",
						 "100111010010100000101010",
						 "100111010010100011011100",
						 "100111010010100110001110",
						 "100111010010101001000000",
						 "100111010001111111010010",
						 "100111010010000010000011",
						 "100111010010000100110100",
						 "100111010010000111100101",
						 "100111010010001010010110",
						 "100111010010001101000111",
						 "100111010010001111111000",
						 "100111010010010010101001",
						 "100111010010010101011010",
						 "100111010010011000001011",
						 "100111010010011010111100",
						 "100111010010011101101101",
						 "100111010010100000011110",
						 "100111010010100011001111",
						 "100111010010100110000000",
						 "100111010010101000110001",
						 "100111010001111111010010",
						 "100111010010000010000011",
						 "100111010010000100110100",
						 "100111010010000111100101",
						 "100111010010001010010110",
						 "100111010010001101000111",
						 "100111010010001111111000",
						 "100111010010010010101001",
						 "100111010010010101011010",
						 "100111010010011000001011",
						 "100111010010011010111100",
						 "100111010010011101101101",
						 "100111010010100000011110",
						 "100111010010100011001111",
						 "100111010010100110000000",
						 "100111010010101000110001",
						 "100111010100100010010000",
						 "100111010100100101000001",
						 "100111010100100111110010",
						 "100111010100101010100011",
						 "100111010100101101010100",
						 "100111010100110000000101",
						 "100111010100110010110110",
						 "100111010100110101100111",
						 "100111010100111000011000",
						 "100111010100111011001001",
						 "100111010100111101111010",
						 "100111010101000000101011",
						 "100111010101000011011100",
						 "100111010101000110001101",
						 "100111010101001000111110",
						 "100111010101001011101111",
						 "100111010100100010010000",
						 "100111010100100101000001",
						 "100111010100100111110010",
						 "100111010100101010100011",
						 "100111010100101101010100",
						 "100111010100110000000101",
						 "100111010100110010110110",
						 "100111010100110101100111",
						 "100111010100111000011000",
						 "100111010100111011001001",
						 "100111010100111101111010",
						 "100111010101000000101011",
						 "100111010101000011011100",
						 "100111010101000110001101",
						 "100111010101001000111110",
						 "100111010101001011101111",
						 "100111010100100010010000",
						 "100111010100100101000000",
						 "100111010100100111110000",
						 "100111010100101010100000",
						 "100111010100101101010000",
						 "100111010100110000000000",
						 "100111010100110010110000",
						 "100111010100110101100000",
						 "100111010100111000010000",
						 "100111010100111011000000",
						 "100111010100111101110000",
						 "100111010101000000100000",
						 "100111010101000011010000",
						 "100111010101000110000000",
						 "100111010101001000110000",
						 "100111010101001011100000",
						 "100111010100100010010000",
						 "100111010100100101000000",
						 "100111010100100111110000",
						 "100111010100101010100000",
						 "100111010100101101010000",
						 "100111010100110000000000",
						 "100111010100110010110000",
						 "100111010100110101100000",
						 "100111010100111000010000",
						 "100111010100111011000000",
						 "100111010100111101110000",
						 "100111010101000000100000",
						 "100111010101000011010000",
						 "100111010101000110000000",
						 "100111010101001000110000",
						 "100111010101001011100000",
						 "100111010111000101001110",
						 "100111010111000111111110",
						 "100111010111001010101110",
						 "100111010111001101011110",
						 "100111010111010000001110",
						 "100111010111010010111110",
						 "100111010111010101101110",
						 "100111010111011000011110",
						 "100111010111011011001110",
						 "100111010111011101111110",
						 "100111010111100000101110",
						 "100111010111100011011110",
						 "100111010111100110001110",
						 "100111010111101000111110",
						 "100111010111101011101110",
						 "100111010111101110011110",
						 "100111010111000101001110",
						 "100111010111000111111101",
						 "100111010111001010101100",
						 "100111010111001101011011",
						 "100111010111010000001010",
						 "100111010111010010111001",
						 "100111010111010101101000",
						 "100111010111011000010111",
						 "100111010111011011000110",
						 "100111010111011101110101",
						 "100111010111100000100100",
						 "100111010111100011010011",
						 "100111010111100110000010",
						 "100111010111101000110001",
						 "100111010111101011100000",
						 "100111010111101110001111",
						 "100111010111000101001110",
						 "100111010111000111111101",
						 "100111010111001010101100",
						 "100111010111001101011011",
						 "100111010111010000001010",
						 "100111010111010010111001",
						 "100111010111010101101000",
						 "100111010111011000010111",
						 "100111010111011011000110",
						 "100111010111011101110101",
						 "100111010111100000100100",
						 "100111010111100011010011",
						 "100111010111100110000010",
						 "100111010111101000110001",
						 "100111010111101011100000",
						 "100111010111101110001111",
						 "100111010111000101001110",
						 "100111010111000111111101",
						 "100111010111001010101100",
						 "100111010111001101011011",
						 "100111010111010000001010",
						 "100111010111010010111001",
						 "100111010111010101101000",
						 "100111010111011000010111",
						 "100111010111011011000110",
						 "100111010111011101110101",
						 "100111010111100000100100",
						 "100111010111100011010011",
						 "100111010111100110000010",
						 "100111010111101000110001",
						 "100111010111101011100000",
						 "100111010111101110001111",
						 "100111011001101000001100",
						 "100111011001101010111011",
						 "100111011001101101101010",
						 "100111011001110000011001",
						 "100111011001110011001000",
						 "100111011001110101110111",
						 "100111011001111000100110",
						 "100111011001111011010101",
						 "100111011001111110000100",
						 "100111011010000000110011",
						 "100111011010000011100010",
						 "100111011010000110010001",
						 "100111011010001001000000",
						 "100111011010001011101111",
						 "100111011010001110011110",
						 "100111011010010001001101",
						 "100111011001101000001100",
						 "100111011001101010111010",
						 "100111011001101101101000",
						 "100111011001110000010110",
						 "100111011001110011000100",
						 "100111011001110101110010",
						 "100111011001111000100000",
						 "100111011001111011001110",
						 "100111011001111101111100",
						 "100111011010000000101010",
						 "100111011010000011011000",
						 "100111011010000110000110",
						 "100111011010001000110100",
						 "100111011010001011100010",
						 "100111011010001110010000",
						 "100111011010010000111110",
						 "100111011001101000001100",
						 "100111011001101010111010",
						 "100111011001101101101000",
						 "100111011001110000010110",
						 "100111011001110011000100",
						 "100111011001110101110010",
						 "100111011001111000100000",
						 "100111011001111011001110",
						 "100111011001111101111100",
						 "100111011010000000101010",
						 "100111011010000011011000",
						 "100111011010000110000110",
						 "100111011010001000110100",
						 "100111011010001011100010",
						 "100111011010001110010000",
						 "100111011010010000111110",
						 "100111011100001011001010",
						 "100111011100001101111000",
						 "100111011100010000100110",
						 "100111011100010011010100",
						 "100111011100010110000010",
						 "100111011100011000110000",
						 "100111011100011011011110",
						 "100111011100011110001100",
						 "100111011100100000111010",
						 "100111011100100011101000",
						 "100111011100100110010110",
						 "100111011100101001000100",
						 "100111011100101011110010",
						 "100111011100101110100000",
						 "100111011100110001001110",
						 "100111011100110011111100",
						 "100111011100001011001010",
						 "100111011100001101110111",
						 "100111011100010000100100",
						 "100111011100010011010001",
						 "100111011100010101111110",
						 "100111011100011000101011",
						 "100111011100011011011000",
						 "100111011100011110000101",
						 "100111011100100000110010",
						 "100111011100100011011111",
						 "100111011100100110001100",
						 "100111011100101000111001",
						 "100111011100101011100110",
						 "100111011100101110010011",
						 "100111011100110001000000",
						 "100111011100110011101101",
						 "100111011100001011001010",
						 "100111011100001101110111",
						 "100111011100010000100100",
						 "100111011100010011010001",
						 "100111011100010101111110",
						 "100111011100011000101011",
						 "100111011100011011011000",
						 "100111011100011110000101",
						 "100111011100100000110010",
						 "100111011100100011011111",
						 "100111011100100110001100",
						 "100111011100101000111001",
						 "100111011100101011100110",
						 "100111011100101110010011",
						 "100111011100110001000000",
						 "100111011100110011101101",
						 "100111011100001011001010",
						 "100111011100001101110111",
						 "100111011100010000100100",
						 "100111011100010011010001",
						 "100111011100010101111110",
						 "100111011100011000101011",
						 "100111011100011011011000",
						 "100111011100011110000101",
						 "100111011100100000110010",
						 "100111011100100011011111",
						 "100111011100100110001100",
						 "100111011100101000111001",
						 "100111011100101011100110",
						 "100111011100101110010011",
						 "100111011100110001000000",
						 "100111011100110011101101",
						 "100111011110101110001000",
						 "100111011110110000110101",
						 "100111011110110011100010",
						 "100111011110110110001111",
						 "100111011110111000111100",
						 "100111011110111011101001",
						 "100111011110111110010110",
						 "100111011111000001000011",
						 "100111011111000011110000",
						 "100111011111000110011101",
						 "100111011111001001001010",
						 "100111011111001011110111",
						 "100111011111001110100100",
						 "100111011111010001010001",
						 "100111011111010011111110",
						 "100111011111010110101011",
						 "100111011110101110001000",
						 "100111011110110000110100",
						 "100111011110110011100000",
						 "100111011110110110001100",
						 "100111011110111000111000",
						 "100111011110111011100100",
						 "100111011110111110010000",
						 "100111011111000000111100",
						 "100111011111000011101000",
						 "100111011111000110010100",
						 "100111011111001001000000",
						 "100111011111001011101100",
						 "100111011111001110011000",
						 "100111011111010001000100",
						 "100111011111010011110000",
						 "100111011111010110011100",
						 "100111011110101110001000",
						 "100111011110110000110100",
						 "100111011110110011100000",
						 "100111011110110110001100",
						 "100111011110111000111000",
						 "100111011110111011100100",
						 "100111011110111110010000",
						 "100111011111000000111100",
						 "100111011111000011101000",
						 "100111011111000110010100",
						 "100111011111001001000000",
						 "100111011111001011101100",
						 "100111011111001110011000",
						 "100111011111010001000100",
						 "100111011111010011110000",
						 "100111011111010110011100",
						 "100111011110101110001000",
						 "100111011110110000110100",
						 "100111011110110011100000",
						 "100111011110110110001100",
						 "100111011110111000111000",
						 "100111011110111011100100",
						 "100111011110111110010000",
						 "100111011111000000111100",
						 "100111011111000011101000",
						 "100111011111000110010100",
						 "100111011111001001000000",
						 "100111011111001011101100",
						 "100111011111001110011000",
						 "100111011111010001000100",
						 "100111011111010011110000",
						 "100111011111010110011100",
						 "100111100001010001000110",
						 "100111100001010011110001",
						 "100111100001010110011100",
						 "100111100001011001000111",
						 "100111100001011011110010",
						 "100111100001011110011101",
						 "100111100001100001001000",
						 "100111100001100011110011",
						 "100111100001100110011110",
						 "100111100001101001001001",
						 "100111100001101011110100",
						 "100111100001101110011111",
						 "100111100001110001001010",
						 "100111100001110011110101",
						 "100111100001110110100000",
						 "100111100001111001001011",
						 "100111100001010001000110",
						 "100111100001010011110001",
						 "100111100001010110011100",
						 "100111100001011001000111",
						 "100111100001011011110010",
						 "100111100001011110011101",
						 "100111100001100001001000",
						 "100111100001100011110011",
						 "100111100001100110011110",
						 "100111100001101001001001",
						 "100111100001101011110100",
						 "100111100001101110011111",
						 "100111100001110001001010",
						 "100111100001110011110101",
						 "100111100001110110100000",
						 "100111100001111001001011",
						 "100111100001010001000110",
						 "100111100001010011110001",
						 "100111100001010110011100",
						 "100111100001011001000111",
						 "100111100001011011110010",
						 "100111100001011110011101",
						 "100111100001100001001000",
						 "100111100001100011110011",
						 "100111100001100110011110",
						 "100111100001101001001001",
						 "100111100001101011110100",
						 "100111100001101110011111",
						 "100111100001110001001010",
						 "100111100001110011110101",
						 "100111100001110110100000",
						 "100111100001111001001011",
						 "100111100001010001000110",
						 "100111100001010011110001",
						 "100111100001010110011100",
						 "100111100001011001000111",
						 "100111100001011011110010",
						 "100111100001011110011101",
						 "100111100001100001001000",
						 "100111100001100011110011",
						 "100111100001100110011110",
						 "100111100001101001001001",
						 "100111100001101011110100",
						 "100111100001101110011111",
						 "100111100001110001001010",
						 "100111100001110011110101",
						 "100111100001110110100000",
						 "100111100001111001001011",
						 "100111100011110100000100",
						 "100111100011110110101110",
						 "100111100011111001011000",
						 "100111100011111100000010",
						 "100111100011111110101100",
						 "100111100100000001010110",
						 "100111100100000100000000",
						 "100111100100000110101010",
						 "100111100100001001010100",
						 "100111100100001011111110",
						 "100111100100001110101000",
						 "100111100100010001010010",
						 "100111100100010011111100",
						 "100111100100010110100110",
						 "100111100100011001010000",
						 "100111100100011011111010",
						 "100111100011110100000100",
						 "100111100011110110101110",
						 "100111100011111001011000",
						 "100111100011111100000010",
						 "100111100011111110101100",
						 "100111100100000001010110",
						 "100111100100000100000000",
						 "100111100100000110101010",
						 "100111100100001001010100",
						 "100111100100001011111110",
						 "100111100100001110101000",
						 "100111100100010001010010",
						 "100111100100010011111100",
						 "100111100100010110100110",
						 "100111100100011001010000",
						 "100111100100011011111010",
						 "100111100011110100000100",
						 "100111100011110110101110",
						 "100111100011111001011000",
						 "100111100011111100000010",
						 "100111100011111110101100",
						 "100111100100000001010110",
						 "100111100100000100000000",
						 "100111100100000110101010",
						 "100111100100001001010100",
						 "100111100100001011111110",
						 "100111100100001110101000",
						 "100111100100010001010010",
						 "100111100100010011111100",
						 "100111100100010110100110",
						 "100111100100011001010000",
						 "100111100100011011111010",
						 "100111100110010111000010",
						 "100111100110011001101011",
						 "100111100110011100010100",
						 "100111100110011110111101",
						 "100111100110100001100110",
						 "100111100110100100001111",
						 "100111100110100110111000",
						 "100111100110101001100001",
						 "100111100110101100001010",
						 "100111100110101110110011",
						 "100111100110110001011100",
						 "100111100110110100000101",
						 "100111100110110110101110",
						 "100111100110111001010111",
						 "100111100110111100000000",
						 "100111100110111110101001",
						 "100111100110010111000010",
						 "100111100110011001101011",
						 "100111100110011100010100",
						 "100111100110011110111101",
						 "100111100110100001100110",
						 "100111100110100100001111",
						 "100111100110100110111000",
						 "100111100110101001100001",
						 "100111100110101100001010",
						 "100111100110101110110011",
						 "100111100110110001011100",
						 "100111100110110100000101",
						 "100111100110110110101110",
						 "100111100110111001010111",
						 "100111100110111100000000",
						 "100111100110111110101001",
						 "100111100110010111000010",
						 "100111100110011001101011",
						 "100111100110011100010100",
						 "100111100110011110111101",
						 "100111100110100001100110",
						 "100111100110100100001111",
						 "100111100110100110111000",
						 "100111100110101001100001",
						 "100111100110101100001010",
						 "100111100110101110110011",
						 "100111100110110001011100",
						 "100111100110110100000101",
						 "100111100110110110101110",
						 "100111100110111001010111",
						 "100111100110111100000000",
						 "100111100110111110101001",
						 "100111100110010111000010",
						 "100111100110011001101010",
						 "100111100110011100010010",
						 "100111100110011110111010",
						 "100111100110100001100010",
						 "100111100110100100001010",
						 "100111100110100110110010",
						 "100111100110101001011010",
						 "100111100110101100000010",
						 "100111100110101110101010",
						 "100111100110110001010010",
						 "100111100110110011111010",
						 "100111100110110110100010",
						 "100111100110111001001010",
						 "100111100110111011110010",
						 "100111100110111110011010",
						 "100111101000111010000000",
						 "100111101000111100101000",
						 "100111101000111111010000",
						 "100111101001000001111000",
						 "100111101001000100100000",
						 "100111101001000111001000",
						 "100111101001001001110000",
						 "100111101001001100011000",
						 "100111101001001111000000",
						 "100111101001010001101000",
						 "100111101001010100010000",
						 "100111101001010110111000",
						 "100111101001011001100000",
						 "100111101001011100001000",
						 "100111101001011110110000",
						 "100111101001100001011000",
						 "100111101000111010000000",
						 "100111101000111100101000",
						 "100111101000111111010000",
						 "100111101001000001111000",
						 "100111101001000100100000",
						 "100111101001000111001000",
						 "100111101001001001110000",
						 "100111101001001100011000",
						 "100111101001001111000000",
						 "100111101001010001101000",
						 "100111101001010100010000",
						 "100111101001010110111000",
						 "100111101001011001100000",
						 "100111101001011100001000",
						 "100111101001011110110000",
						 "100111101001100001011000",
						 "100111101000111010000000",
						 "100111101000111100101000",
						 "100111101000111111010000",
						 "100111101001000001111000",
						 "100111101001000100100000",
						 "100111101001000111001000",
						 "100111101001001001110000",
						 "100111101001001100011000",
						 "100111101001001111000000",
						 "100111101001010001101000",
						 "100111101001010100010000",
						 "100111101001010110111000",
						 "100111101001011001100000",
						 "100111101001011100001000",
						 "100111101001011110110000",
						 "100111101001100001011000",
						 "100111101000111010000000",
						 "100111101000111100100111",
						 "100111101000111111001110",
						 "100111101001000001110101",
						 "100111101001000100011100",
						 "100111101001000111000011",
						 "100111101001001001101010",
						 "100111101001001100010001",
						 "100111101001001110111000",
						 "100111101001010001011111",
						 "100111101001010100000110",
						 "100111101001010110101101",
						 "100111101001011001010100",
						 "100111101001011011111011",
						 "100111101001011110100010",
						 "100111101001100001001001",
						 "100111101011011100111110",
						 "100111101011011111100101",
						 "100111101011100010001100",
						 "100111101011100100110011",
						 "100111101011100111011010",
						 "100111101011101010000001",
						 "100111101011101100101000",
						 "100111101011101111001111",
						 "100111101011110001110110",
						 "100111101011110100011101",
						 "100111101011110111000100",
						 "100111101011111001101011",
						 "100111101011111100010010",
						 "100111101011111110111001",
						 "100111101100000001100000",
						 "100111101100000100000111",
						 "100111101011011100111110",
						 "100111101011011111100101",
						 "100111101011100010001100",
						 "100111101011100100110011",
						 "100111101011100111011010",
						 "100111101011101010000001",
						 "100111101011101100101000",
						 "100111101011101111001111",
						 "100111101011110001110110",
						 "100111101011110100011101",
						 "100111101011110111000100",
						 "100111101011111001101011",
						 "100111101011111100010010",
						 "100111101011111110111001",
						 "100111101100000001100000",
						 "100111101100000100000111",
						 "100111101011011100111110",
						 "100111101011011111100100",
						 "100111101011100010001010",
						 "100111101011100100110000",
						 "100111101011100111010110",
						 "100111101011101001111100",
						 "100111101011101100100010",
						 "100111101011101111001000",
						 "100111101011110001101110",
						 "100111101011110100010100",
						 "100111101011110110111010",
						 "100111101011111001100000",
						 "100111101011111100000110",
						 "100111101011111110101100",
						 "100111101100000001010010",
						 "100111101100000011111000",
						 "100111101011011100111110",
						 "100111101011011111100100",
						 "100111101011100010001010",
						 "100111101011100100110000",
						 "100111101011100111010110",
						 "100111101011101001111100",
						 "100111101011101100100010",
						 "100111101011101111001000",
						 "100111101011110001101110",
						 "100111101011110100010100",
						 "100111101011110110111010",
						 "100111101011111001100000",
						 "100111101011111100000110",
						 "100111101011111110101100",
						 "100111101100000001010010",
						 "100111101100000011111000",
						 "100111101101111111111100",
						 "100111101110000010100010",
						 "100111101110000101001000",
						 "100111101110000111101110",
						 "100111101110001010010100",
						 "100111101110001100111010",
						 "100111101110001111100000",
						 "100111101110010010000110",
						 "100111101110010100101100",
						 "100111101110010111010010",
						 "100111101110011001111000",
						 "100111101110011100011110",
						 "100111101110011111000100",
						 "100111101110100001101010",
						 "100111101110100100010000",
						 "100111101110100110110110",
						 "100111101101111111111100",
						 "100111101110000010100010",
						 "100111101110000101001000",
						 "100111101110000111101110",
						 "100111101110001010010100",
						 "100111101110001100111010",
						 "100111101110001111100000",
						 "100111101110010010000110",
						 "100111101110010100101100",
						 "100111101110010111010010",
						 "100111101110011001111000",
						 "100111101110011100011110",
						 "100111101110011111000100",
						 "100111101110100001101010",
						 "100111101110100100010000",
						 "100111101110100110110110",
						 "100111101101111111111100",
						 "100111101110000010100001",
						 "100111101110000101000110",
						 "100111101110000111101011",
						 "100111101110001010010000",
						 "100111101110001100110101",
						 "100111101110001111011010",
						 "100111101110010001111111",
						 "100111101110010100100100",
						 "100111101110010111001001",
						 "100111101110011001101110",
						 "100111101110011100010011",
						 "100111101110011110111000",
						 "100111101110100001011101",
						 "100111101110100100000010",
						 "100111101110100110100111",
						 "100111101101111111111100",
						 "100111101110000010100001",
						 "100111101110000101000110",
						 "100111101110000111101011",
						 "100111101110001010010000",
						 "100111101110001100110101",
						 "100111101110001111011010",
						 "100111101110010001111111",
						 "100111101110010100100100",
						 "100111101110010111001001",
						 "100111101110011001101110",
						 "100111101110011100010011",
						 "100111101110011110111000",
						 "100111101110100001011101",
						 "100111101110100100000010",
						 "100111101110100110100111",
						 "100111110000100010111010",
						 "100111110000100101011111",
						 "100111110000101000000100",
						 "100111110000101010101001",
						 "100111110000101101001110",
						 "100111110000101111110011",
						 "100111110000110010011000",
						 "100111110000110100111101",
						 "100111110000110111100010",
						 "100111110000111010000111",
						 "100111110000111100101100",
						 "100111110000111111010001",
						 "100111110001000001110110",
						 "100111110001000100011011",
						 "100111110001000111000000",
						 "100111110001001001100101",
						 "100111110000100010111010",
						 "100111110000100101011110",
						 "100111110000101000000010",
						 "100111110000101010100110",
						 "100111110000101101001010",
						 "100111110000101111101110",
						 "100111110000110010010010",
						 "100111110000110100110110",
						 "100111110000110111011010",
						 "100111110000111001111110",
						 "100111110000111100100010",
						 "100111110000111111000110",
						 "100111110001000001101010",
						 "100111110001000100001110",
						 "100111110001000110110010",
						 "100111110001001001010110",
						 "100111110000100010111010",
						 "100111110000100101011110",
						 "100111110000101000000010",
						 "100111110000101010100110",
						 "100111110000101101001010",
						 "100111110000101111101110",
						 "100111110000110010010010",
						 "100111110000110100110110",
						 "100111110000110111011010",
						 "100111110000111001111110",
						 "100111110000111100100010",
						 "100111110000111111000110",
						 "100111110001000001101010",
						 "100111110001000100001110",
						 "100111110001000110110010",
						 "100111110001001001010110",
						 "100111110000100010111010",
						 "100111110000100101011110",
						 "100111110000101000000010",
						 "100111110000101010100110",
						 "100111110000101101001010",
						 "100111110000101111101110",
						 "100111110000110010010010",
						 "100111110000110100110110",
						 "100111110000110111011010",
						 "100111110000111001111110",
						 "100111110000111100100010",
						 "100111110000111111000110",
						 "100111110001000001101010",
						 "100111110001000100001110",
						 "100111110001000110110010",
						 "100111110001001001010110",
						 "100111110011000101111000",
						 "100111110011001000011011",
						 "100111110011001010111110",
						 "100111110011001101100001",
						 "100111110011010000000100",
						 "100111110011010010100111",
						 "100111110011010101001010",
						 "100111110011010111101101",
						 "100111110011011010010000",
						 "100111110011011100110011",
						 "100111110011011111010110",
						 "100111110011100001111001",
						 "100111110011100100011100",
						 "100111110011100110111111",
						 "100111110011101001100010",
						 "100111110011101100000101",
						 "100111110011000101111000",
						 "100111110011001000011011",
						 "100111110011001010111110",
						 "100111110011001101100001",
						 "100111110011010000000100",
						 "100111110011010010100111",
						 "100111110011010101001010",
						 "100111110011010111101101",
						 "100111110011011010010000",
						 "100111110011011100110011",
						 "100111110011011111010110",
						 "100111110011100001111001",
						 "100111110011100100011100",
						 "100111110011100110111111",
						 "100111110011101001100010",
						 "100111110011101100000101",
						 "100111110011000101111000",
						 "100111110011001000011011",
						 "100111110011001010111110",
						 "100111110011001101100001",
						 "100111110011010000000100",
						 "100111110011010010100111",
						 "100111110011010101001010",
						 "100111110011010111101101",
						 "100111110011011010010000",
						 "100111110011011100110011",
						 "100111110011011111010110",
						 "100111110011100001111001",
						 "100111110011100100011100",
						 "100111110011100110111111",
						 "100111110011101001100010",
						 "100111110011101100000101",
						 "100111110011000101111000",
						 "100111110011001000011011",
						 "100111110011001010111110",
						 "100111110011001101100001",
						 "100111110011010000000100",
						 "100111110011010010100111",
						 "100111110011010101001010",
						 "100111110011010111101101",
						 "100111110011011010010000",
						 "100111110011011100110011",
						 "100111110011011111010110",
						 "100111110011100001111001",
						 "100111110011100100011100",
						 "100111110011100110111111",
						 "100111110011101001100010",
						 "100111110011101100000101",
						 "100111110101101000110110",
						 "100111110101101011011000",
						 "100111110101101101111010",
						 "100111110101110000011100",
						 "100111110101110010111110",
						 "100111110101110101100000",
						 "100111110101111000000010",
						 "100111110101111010100100",
						 "100111110101111101000110",
						 "100111110101111111101000",
						 "100111110110000010001010",
						 "100111110110000100101100",
						 "100111110110000111001110",
						 "100111110110001001110000",
						 "100111110110001100010010",
						 "100111110110001110110100",
						 "100111110101101000110110",
						 "100111110101101011011000",
						 "100111110101101101111010",
						 "100111110101110000011100",
						 "100111110101110010111110",
						 "100111110101110101100000",
						 "100111110101111000000010",
						 "100111110101111010100100",
						 "100111110101111101000110",
						 "100111110101111111101000",
						 "100111110110000010001010",
						 "100111110110000100101100",
						 "100111110110000111001110",
						 "100111110110001001110000",
						 "100111110110001100010010",
						 "100111110110001110110100",
						 "100111110101101000110110",
						 "100111110101101011011000",
						 "100111110101101101111010",
						 "100111110101110000011100",
						 "100111110101110010111110",
						 "100111110101110101100000",
						 "100111110101111000000010",
						 "100111110101111010100100",
						 "100111110101111101000110",
						 "100111110101111111101000",
						 "100111110110000010001010",
						 "100111110110000100101100",
						 "100111110110000111001110",
						 "100111110110001001110000",
						 "100111110110001100010010",
						 "100111110110001110110100",
						 "100111110101101000110110",
						 "100111110101101011010111",
						 "100111110101101101111000",
						 "100111110101110000011001",
						 "100111110101110010111010",
						 "100111110101110101011011",
						 "100111110101110111111100",
						 "100111110101111010011101",
						 "100111110101111100111110",
						 "100111110101111111011111",
						 "100111110110000010000000",
						 "100111110110000100100001",
						 "100111110110000111000010",
						 "100111110110001001100011",
						 "100111110110001100000100",
						 "100111110110001110100101",
						 "100111111000001011110100",
						 "100111111000001110010101",
						 "100111111000010000110110",
						 "100111111000010011010111",
						 "100111111000010101111000",
						 "100111111000011000011001",
						 "100111111000011010111010",
						 "100111111000011101011011",
						 "100111111000011111111100",
						 "100111111000100010011101",
						 "100111111000100100111110",
						 "100111111000100111011111",
						 "100111111000101010000000",
						 "100111111000101100100001",
						 "100111111000101111000010",
						 "100111111000110001100011",
						 "100111111000001011110100",
						 "100111111000001110010101",
						 "100111111000010000110110",
						 "100111111000010011010111",
						 "100111111000010101111000",
						 "100111111000011000011001",
						 "100111111000011010111010",
						 "100111111000011101011011",
						 "100111111000011111111100",
						 "100111111000100010011101",
						 "100111111000100100111110",
						 "100111111000100111011111",
						 "100111111000101010000000",
						 "100111111000101100100001",
						 "100111111000101111000010",
						 "100111111000110001100011",
						 "100111111000001011110100",
						 "100111111000001110010100",
						 "100111111000010000110100",
						 "100111111000010011010100",
						 "100111111000010101110100",
						 "100111111000011000010100",
						 "100111111000011010110100",
						 "100111111000011101010100",
						 "100111111000011111110100",
						 "100111111000100010010100",
						 "100111111000100100110100",
						 "100111111000100111010100",
						 "100111111000101001110100",
						 "100111111000101100010100",
						 "100111111000101110110100",
						 "100111111000110001010100",
						 "100111111000001011110100",
						 "100111111000001110010100",
						 "100111111000010000110100",
						 "100111111000010011010100",
						 "100111111000010101110100",
						 "100111111000011000010100",
						 "100111111000011010110100",
						 "100111111000011101010100",
						 "100111111000011111110100",
						 "100111111000100010010100",
						 "100111111000100100110100",
						 "100111111000100111010100",
						 "100111111000101001110100",
						 "100111111000101100010100",
						 "100111111000101110110100",
						 "100111111000110001010100",
						 "100111111010101110110010",
						 "100111111010110001010010",
						 "100111111010110011110010",
						 "100111111010110110010010",
						 "100111111010111000110010",
						 "100111111010111011010010",
						 "100111111010111101110010",
						 "100111111011000000010010",
						 "100111111011000010110010",
						 "100111111011000101010010",
						 "100111111011000111110010",
						 "100111111011001010010010",
						 "100111111011001100110010",
						 "100111111011001111010010",
						 "100111111011010001110010",
						 "100111111011010100010010",
						 "100111111010101110110010",
						 "100111111010110001010001",
						 "100111111010110011110000",
						 "100111111010110110001111",
						 "100111111010111000101110",
						 "100111111010111011001101",
						 "100111111010111101101100",
						 "100111111011000000001011",
						 "100111111011000010101010",
						 "100111111011000101001001",
						 "100111111011000111101000",
						 "100111111011001010000111",
						 "100111111011001100100110",
						 "100111111011001111000101",
						 "100111111011010001100100",
						 "100111111011010100000011",
						 "100111111010101110110010",
						 "100111111010110001010001",
						 "100111111010110011110000",
						 "100111111010110110001111",
						 "100111111010111000101110",
						 "100111111010111011001101",
						 "100111111010111101101100",
						 "100111111011000000001011",
						 "100111111011000010101010",
						 "100111111011000101001001",
						 "100111111011000111101000",
						 "100111111011001010000111",
						 "100111111011001100100110",
						 "100111111011001111000101",
						 "100111111011010001100100",
						 "100111111011010100000011",
						 "100111111010101110110010",
						 "100111111010110001010001",
						 "100111111010110011110000",
						 "100111111010110110001111",
						 "100111111010111000101110",
						 "100111111010111011001101",
						 "100111111010111101101100",
						 "100111111011000000001011",
						 "100111111011000010101010",
						 "100111111011000101001001",
						 "100111111011000111101000",
						 "100111111011001010000111",
						 "100111111011001100100110",
						 "100111111011001111000101",
						 "100111111011010001100100",
						 "100111111011010100000011",
						 "100111111101010001110000",
						 "100111111101010100001111",
						 "100111111101010110101110",
						 "100111111101011001001101",
						 "100111111101011011101100",
						 "100111111101011110001011",
						 "100111111101100000101010",
						 "100111111101100011001001",
						 "100111111101100101101000",
						 "100111111101101000000111",
						 "100111111101101010100110",
						 "100111111101101101000101",
						 "100111111101101111100100",
						 "100111111101110010000011",
						 "100111111101110100100010",
						 "100111111101110111000001",
						 "100111111101010001110000",
						 "100111111101010100001110",
						 "100111111101010110101100",
						 "100111111101011001001010",
						 "100111111101011011101000",
						 "100111111101011110000110",
						 "100111111101100000100100",
						 "100111111101100011000010",
						 "100111111101100101100000",
						 "100111111101100111111110",
						 "100111111101101010011100",
						 "100111111101101100111010",
						 "100111111101101111011000",
						 "100111111101110001110110",
						 "100111111101110100010100",
						 "100111111101110110110010",
						 "100111111101010001110000",
						 "100111111101010100001110",
						 "100111111101010110101100",
						 "100111111101011001001010",
						 "100111111101011011101000",
						 "100111111101011110000110",
						 "100111111101100000100100",
						 "100111111101100011000010",
						 "100111111101100101100000",
						 "100111111101100111111110",
						 "100111111101101010011100",
						 "100111111101101100111010",
						 "100111111101101111011000",
						 "100111111101110001110110",
						 "100111111101110100010100",
						 "100111111101110110110010",
						 "100111111101010001110000",
						 "100111111101010100001110",
						 "100111111101010110101100",
						 "100111111101011001001010",
						 "100111111101011011101000",
						 "100111111101011110000110",
						 "100111111101100000100100",
						 "100111111101100011000010",
						 "100111111101100101100000",
						 "100111111101100111111110",
						 "100111111101101010011100",
						 "100111111101101100111010",
						 "100111111101101111011000",
						 "100111111101110001110110",
						 "100111111101110100010100",
						 "100111111101110110110010",
						 "100111111111110100101110",
						 "100111111111110111001011",
						 "100111111111111001101000",
						 "100111111111111100000101",
						 "100111111111111110100010",
						 "101000000000000000111111",
						 "101000000000000011011100",
						 "101000000000000101111001",
						 "101000000000001000010110",
						 "101000000000001010110011",
						 "101000000000001101010000",
						 "101000000000001111101101",
						 "101000000000010010001010",
						 "101000000000010100100111",
						 "101000000000010111000100",
						 "101000000000011001100001",
						 "100111111111110100101110",
						 "100111111111110111001011",
						 "100111111111111001101000",
						 "100111111111111100000101",
						 "100111111111111110100010",
						 "101000000000000000111111",
						 "101000000000000011011100",
						 "101000000000000101111001",
						 "101000000000001000010110",
						 "101000000000001010110011",
						 "101000000000001101010000",
						 "101000000000001111101101",
						 "101000000000010010001010",
						 "101000000000010100100111",
						 "101000000000010111000100",
						 "101000000000011001100001",
						 "100111111111110100101110",
						 "100111111111110111001011",
						 "100111111111111001101000",
						 "100111111111111100000101",
						 "100111111111111110100010",
						 "101000000000000000111111",
						 "101000000000000011011100",
						 "101000000000000101111001",
						 "101000000000001000010110",
						 "101000000000001010110011",
						 "101000000000001101010000",
						 "101000000000001111101101",
						 "101000000000010010001010",
						 "101000000000010100100111",
						 "101000000000010111000100",
						 "101000000000011001100001",
						 "100111111111110100101110",
						 "100111111111110111001010",
						 "100111111111111001100110",
						 "100111111111111100000010",
						 "100111111111111110011110",
						 "101000000000000000111010",
						 "101000000000000011010110",
						 "101000000000000101110010",
						 "101000000000001000001110",
						 "101000000000001010101010",
						 "101000000000001101000110",
						 "101000000000001111100010",
						 "101000000000010001111110",
						 "101000000000010100011010",
						 "101000000000010110110110",
						 "101000000000011001010010",
						 "101000000010010111101100",
						 "101000000010011010001000",
						 "101000000010011100100100",
						 "101000000010011111000000",
						 "101000000010100001011100",
						 "101000000010100011111000",
						 "101000000010100110010100",
						 "101000000010101000110000",
						 "101000000010101011001100",
						 "101000000010101101101000",
						 "101000000010110000000100",
						 "101000000010110010100000",
						 "101000000010110100111100",
						 "101000000010110111011000",
						 "101000000010111001110100",
						 "101000000010111100010000",
						 "101000000010010111101100",
						 "101000000010011010001000",
						 "101000000010011100100100",
						 "101000000010011111000000",
						 "101000000010100001011100",
						 "101000000010100011111000",
						 "101000000010100110010100",
						 "101000000010101000110000",
						 "101000000010101011001100",
						 "101000000010101101101000",
						 "101000000010110000000100",
						 "101000000010110010100000",
						 "101000000010110100111100",
						 "101000000010110111011000",
						 "101000000010111001110100",
						 "101000000010111100010000",
						 "101000000010010111101100",
						 "101000000010011010000111",
						 "101000000010011100100010",
						 "101000000010011110111101",
						 "101000000010100001011000",
						 "101000000010100011110011",
						 "101000000010100110001110",
						 "101000000010101000101001",
						 "101000000010101011000100",
						 "101000000010101101011111",
						 "101000000010101111111010",
						 "101000000010110010010101",
						 "101000000010110100110000",
						 "101000000010110111001011",
						 "101000000010111001100110",
						 "101000000010111100000001",
						 "101000000010010111101100",
						 "101000000010011010000111",
						 "101000000010011100100010",
						 "101000000010011110111101",
						 "101000000010100001011000",
						 "101000000010100011110011",
						 "101000000010100110001110",
						 "101000000010101000101001",
						 "101000000010101011000100",
						 "101000000010101101011111",
						 "101000000010101111111010",
						 "101000000010110010010101",
						 "101000000010110100110000",
						 "101000000010110111001011",
						 "101000000010111001100110",
						 "101000000010111100000001",
						 "101000000010010111101100",
						 "101000000010011010000111",
						 "101000000010011100100010",
						 "101000000010011110111101",
						 "101000000010100001011000",
						 "101000000010100011110011",
						 "101000000010100110001110",
						 "101000000010101000101001",
						 "101000000010101011000100",
						 "101000000010101101011111",
						 "101000000010101111111010",
						 "101000000010110010010101",
						 "101000000010110100110000",
						 "101000000010110111001011",
						 "101000000010111001100110",
						 "101000000010111100000001",
						 "101000000100111010101010",
						 "101000000100111101000101",
						 "101000000100111111100000",
						 "101000000101000001111011",
						 "101000000101000100010110",
						 "101000000101000110110001",
						 "101000000101001001001100",
						 "101000000101001011100111",
						 "101000000101001110000010",
						 "101000000101010000011101",
						 "101000000101010010111000",
						 "101000000101010101010011",
						 "101000000101010111101110",
						 "101000000101011010001001",
						 "101000000101011100100100",
						 "101000000101011110111111",
						 "101000000100111010101010",
						 "101000000100111101000100",
						 "101000000100111111011110",
						 "101000000101000001111000",
						 "101000000101000100010010",
						 "101000000101000110101100",
						 "101000000101001001000110",
						 "101000000101001011100000",
						 "101000000101001101111010",
						 "101000000101010000010100",
						 "101000000101010010101110",
						 "101000000101010101001000",
						 "101000000101010111100010",
						 "101000000101011001111100",
						 "101000000101011100010110",
						 "101000000101011110110000",
						 "101000000100111010101010",
						 "101000000100111101000100",
						 "101000000100111111011110",
						 "101000000101000001111000",
						 "101000000101000100010010",
						 "101000000101000110101100",
						 "101000000101001001000110",
						 "101000000101001011100000",
						 "101000000101001101111010",
						 "101000000101010000010100",
						 "101000000101010010101110",
						 "101000000101010101001000",
						 "101000000101010111100010",
						 "101000000101011001111100",
						 "101000000101011100010110",
						 "101000000101011110110000",
						 "101000000100111010101010",
						 "101000000100111101000100",
						 "101000000100111111011110",
						 "101000000101000001111000",
						 "101000000101000100010010",
						 "101000000101000110101100",
						 "101000000101001001000110",
						 "101000000101001011100000",
						 "101000000101001101111010",
						 "101000000101010000010100",
						 "101000000101010010101110",
						 "101000000101010101001000",
						 "101000000101010111100010",
						 "101000000101011001111100",
						 "101000000101011100010110",
						 "101000000101011110110000",
						 "101000000111011101101000",
						 "101000000111100000000001",
						 "101000000111100010011010",
						 "101000000111100100110011",
						 "101000000111100111001100",
						 "101000000111101001100101",
						 "101000000111101011111110",
						 "101000000111101110010111",
						 "101000000111110000110000",
						 "101000000111110011001001",
						 "101000000111110101100010",
						 "101000000111110111111011",
						 "101000000111111010010100",
						 "101000000111111100101101",
						 "101000000111111111000110",
						 "101000001000000001011111",
						 "101000000111011101101000",
						 "101000000111100000000001",
						 "101000000111100010011010",
						 "101000000111100100110011",
						 "101000000111100111001100",
						 "101000000111101001100101",
						 "101000000111101011111110",
						 "101000000111101110010111",
						 "101000000111110000110000",
						 "101000000111110011001001",
						 "101000000111110101100010",
						 "101000000111110111111011",
						 "101000000111111010010100",
						 "101000000111111100101101",
						 "101000000111111111000110",
						 "101000001000000001011111",
						 "101000000111011101101000",
						 "101000000111100000000001",
						 "101000000111100010011010",
						 "101000000111100100110011",
						 "101000000111100111001100",
						 "101000000111101001100101",
						 "101000000111101011111110",
						 "101000000111101110010111",
						 "101000000111110000110000",
						 "101000000111110011001001",
						 "101000000111110101100010",
						 "101000000111110111111011",
						 "101000000111111010010100",
						 "101000000111111100101101",
						 "101000000111111111000110",
						 "101000001000000001011111",
						 "101000000111011101101000",
						 "101000000111100000000000",
						 "101000000111100010011000",
						 "101000000111100100110000",
						 "101000000111100111001000",
						 "101000000111101001100000",
						 "101000000111101011111000",
						 "101000000111101110010000",
						 "101000000111110000101000",
						 "101000000111110011000000",
						 "101000000111110101011000",
						 "101000000111110111110000",
						 "101000000111111010001000",
						 "101000000111111100100000",
						 "101000000111111110111000",
						 "101000001000000001010000",
						 "101000001010000000100110",
						 "101000001010000010111110",
						 "101000001010000101010110",
						 "101000001010000111101110",
						 "101000001010001010000110",
						 "101000001010001100011110",
						 "101000001010001110110110",
						 "101000001010010001001110",
						 "101000001010010011100110",
						 "101000001010010101111110",
						 "101000001010011000010110",
						 "101000001010011010101110",
						 "101000001010011101000110",
						 "101000001010011111011110",
						 "101000001010100001110110",
						 "101000001010100100001110",
						 "101000001010000000100110",
						 "101000001010000010111110",
						 "101000001010000101010110",
						 "101000001010000111101110",
						 "101000001010001010000110",
						 "101000001010001100011110",
						 "101000001010001110110110",
						 "101000001010010001001110",
						 "101000001010010011100110",
						 "101000001010010101111110",
						 "101000001010011000010110",
						 "101000001010011010101110",
						 "101000001010011101000110",
						 "101000001010011111011110",
						 "101000001010100001110110",
						 "101000001010100100001110",
						 "101000001010000000100110",
						 "101000001010000010111101",
						 "101000001010000101010100",
						 "101000001010000111101011",
						 "101000001010001010000010",
						 "101000001010001100011001",
						 "101000001010001110110000",
						 "101000001010010001000111",
						 "101000001010010011011110",
						 "101000001010010101110101",
						 "101000001010011000001100",
						 "101000001010011010100011",
						 "101000001010011100111010",
						 "101000001010011111010001",
						 "101000001010100001101000",
						 "101000001010100011111111",
						 "101000001010000000100110",
						 "101000001010000010111101",
						 "101000001010000101010100",
						 "101000001010000111101011",
						 "101000001010001010000010",
						 "101000001010001100011001",
						 "101000001010001110110000",
						 "101000001010010001000111",
						 "101000001010010011011110",
						 "101000001010010101110101",
						 "101000001010011000001100",
						 "101000001010011010100011",
						 "101000001010011100111010",
						 "101000001010011111010001",
						 "101000001010100001101000",
						 "101000001010100011111111",
						 "101000001100100011100100",
						 "101000001100100101111011",
						 "101000001100101000010010",
						 "101000001100101010101001",
						 "101000001100101101000000",
						 "101000001100101111010111",
						 "101000001100110001101110",
						 "101000001100110100000101",
						 "101000001100110110011100",
						 "101000001100111000110011",
						 "101000001100111011001010",
						 "101000001100111101100001",
						 "101000001100111111111000",
						 "101000001101000010001111",
						 "101000001101000100100110",
						 "101000001101000110111101",
						 "101000001100100011100100",
						 "101000001100100101111010",
						 "101000001100101000010000",
						 "101000001100101010100110",
						 "101000001100101100111100",
						 "101000001100101111010010",
						 "101000001100110001101000",
						 "101000001100110011111110",
						 "101000001100110110010100",
						 "101000001100111000101010",
						 "101000001100111011000000",
						 "101000001100111101010110",
						 "101000001100111111101100",
						 "101000001101000010000010",
						 "101000001101000100011000",
						 "101000001101000110101110",
						 "101000001100100011100100",
						 "101000001100100101111010",
						 "101000001100101000010000",
						 "101000001100101010100110",
						 "101000001100101100111100",
						 "101000001100101111010010",
						 "101000001100110001101000",
						 "101000001100110011111110",
						 "101000001100110110010100",
						 "101000001100111000101010",
						 "101000001100111011000000",
						 "101000001100111101010110",
						 "101000001100111111101100",
						 "101000001101000010000010",
						 "101000001101000100011000",
						 "101000001101000110101110",
						 "101000001100100011100100",
						 "101000001100100101111010",
						 "101000001100101000010000",
						 "101000001100101010100110",
						 "101000001100101100111100",
						 "101000001100101111010010",
						 "101000001100110001101000",
						 "101000001100110011111110",
						 "101000001100110110010100",
						 "101000001100111000101010",
						 "101000001100111011000000",
						 "101000001100111101010110",
						 "101000001100111111101100",
						 "101000001101000010000010",
						 "101000001101000100011000",
						 "101000001101000110101110",
						 "101000001100100011100100",
						 "101000001100100101111010",
						 "101000001100101000010000",
						 "101000001100101010100110",
						 "101000001100101100111100",
						 "101000001100101111010010",
						 "101000001100110001101000",
						 "101000001100110011111110",
						 "101000001100110110010100",
						 "101000001100111000101010",
						 "101000001100111011000000",
						 "101000001100111101010110",
						 "101000001100111111101100",
						 "101000001101000010000010",
						 "101000001101000100011000",
						 "101000001101000110101110",
						 "101000001111000110100010",
						 "101000001111001000110111",
						 "101000001111001011001100",
						 "101000001111001101100001",
						 "101000001111001111110110",
						 "101000001111010010001011",
						 "101000001111010100100000",
						 "101000001111010110110101",
						 "101000001111011001001010",
						 "101000001111011011011111",
						 "101000001111011101110100",
						 "101000001111100000001001",
						 "101000001111100010011110",
						 "101000001111100100110011",
						 "101000001111100111001000",
						 "101000001111101001011101",
						 "101000001111000110100010",
						 "101000001111001000110111",
						 "101000001111001011001100",
						 "101000001111001101100001",
						 "101000001111001111110110",
						 "101000001111010010001011",
						 "101000001111010100100000",
						 "101000001111010110110101",
						 "101000001111011001001010",
						 "101000001111011011011111",
						 "101000001111011101110100",
						 "101000001111100000001001",
						 "101000001111100010011110",
						 "101000001111100100110011",
						 "101000001111100111001000",
						 "101000001111101001011101",
						 "101000001111000110100010",
						 "101000001111001000110111",
						 "101000001111001011001100",
						 "101000001111001101100001",
						 "101000001111001111110110",
						 "101000001111010010001011",
						 "101000001111010100100000",
						 "101000001111010110110101",
						 "101000001111011001001010",
						 "101000001111011011011111",
						 "101000001111011101110100",
						 "101000001111100000001001",
						 "101000001111100010011110",
						 "101000001111100100110011",
						 "101000001111100111001000",
						 "101000001111101001011101",
						 "101000001111000110100010",
						 "101000001111001000110110",
						 "101000001111001011001010",
						 "101000001111001101011110",
						 "101000001111001111110010",
						 "101000001111010010000110",
						 "101000001111010100011010",
						 "101000001111010110101110",
						 "101000001111011001000010",
						 "101000001111011011010110",
						 "101000001111011101101010",
						 "101000001111011111111110",
						 "101000001111100010010010",
						 "101000001111100100100110",
						 "101000001111100110111010",
						 "101000001111101001001110",
						 "101000010001101001100000",
						 "101000010001101011110100",
						 "101000010001101110001000",
						 "101000010001110000011100",
						 "101000010001110010110000",
						 "101000010001110101000100",
						 "101000010001110111011000",
						 "101000010001111001101100",
						 "101000010001111100000000",
						 "101000010001111110010100",
						 "101000010010000000101000",
						 "101000010010000010111100",
						 "101000010010000101010000",
						 "101000010010000111100100",
						 "101000010010001001111000",
						 "101000010010001100001100",
						 "101000010001101001100000",
						 "101000010001101011110100",
						 "101000010001101110001000",
						 "101000010001110000011100",
						 "101000010001110010110000",
						 "101000010001110101000100",
						 "101000010001110111011000",
						 "101000010001111001101100",
						 "101000010001111100000000",
						 "101000010001111110010100",
						 "101000010010000000101000",
						 "101000010010000010111100",
						 "101000010010000101010000",
						 "101000010010000111100100",
						 "101000010010001001111000",
						 "101000010010001100001100",
						 "101000010001101001100000",
						 "101000010001101011110011",
						 "101000010001101110000110",
						 "101000010001110000011001",
						 "101000010001110010101100",
						 "101000010001110100111111",
						 "101000010001110111010010",
						 "101000010001111001100101",
						 "101000010001111011111000",
						 "101000010001111110001011",
						 "101000010010000000011110",
						 "101000010010000010110001",
						 "101000010010000101000100",
						 "101000010010000111010111",
						 "101000010010001001101010",
						 "101000010010001011111101",
						 "101000010001101001100000",
						 "101000010001101011110011",
						 "101000010001101110000110",
						 "101000010001110000011001",
						 "101000010001110010101100",
						 "101000010001110100111111",
						 "101000010001110111010010",
						 "101000010001111001100101",
						 "101000010001111011111000",
						 "101000010001111110001011",
						 "101000010010000000011110",
						 "101000010010000010110001",
						 "101000010010000101000100",
						 "101000010010000111010111",
						 "101000010010001001101010",
						 "101000010010001011111101",
						 "101000010001101001100000",
						 "101000010001101011110011",
						 "101000010001101110000110",
						 "101000010001110000011001",
						 "101000010001110010101100",
						 "101000010001110100111111",
						 "101000010001110111010010",
						 "101000010001111001100101",
						 "101000010001111011111000",
						 "101000010001111110001011",
						 "101000010010000000011110",
						 "101000010010000010110001",
						 "101000010010000101000100",
						 "101000010010000111010111",
						 "101000010010001001101010",
						 "101000010010001011111101",
						 "101000010100001100011110",
						 "101000010100001110110000",
						 "101000010100010001000010",
						 "101000010100010011010100",
						 "101000010100010101100110",
						 "101000010100010111111000",
						 "101000010100011010001010",
						 "101000010100011100011100",
						 "101000010100011110101110",
						 "101000010100100001000000",
						 "101000010100100011010010",
						 "101000010100100101100100",
						 "101000010100100111110110",
						 "101000010100101010001000",
						 "101000010100101100011010",
						 "101000010100101110101100",
						 "101000010100001100011110",
						 "101000010100001110110000",
						 "101000010100010001000010",
						 "101000010100010011010100",
						 "101000010100010101100110",
						 "101000010100010111111000",
						 "101000010100011010001010",
						 "101000010100011100011100",
						 "101000010100011110101110",
						 "101000010100100001000000",
						 "101000010100100011010010",
						 "101000010100100101100100",
						 "101000010100100111110110",
						 "101000010100101010001000",
						 "101000010100101100011010",
						 "101000010100101110101100",
						 "101000010100001100011110",
						 "101000010100001110110000",
						 "101000010100010001000010",
						 "101000010100010011010100",
						 "101000010100010101100110",
						 "101000010100010111111000",
						 "101000010100011010001010",
						 "101000010100011100011100",
						 "101000010100011110101110",
						 "101000010100100001000000",
						 "101000010100100011010010",
						 "101000010100100101100100",
						 "101000010100100111110110",
						 "101000010100101010001000",
						 "101000010100101100011010",
						 "101000010100101110101100",
						 "101000010100001100011110",
						 "101000010100001110101111",
						 "101000010100010001000000",
						 "101000010100010011010001",
						 "101000010100010101100010",
						 "101000010100010111110011",
						 "101000010100011010000100",
						 "101000010100011100010101",
						 "101000010100011110100110",
						 "101000010100100000110111",
						 "101000010100100011001000",
						 "101000010100100101011001",
						 "101000010100100111101010",
						 "101000010100101001111011",
						 "101000010100101100001100",
						 "101000010100101110011101",
						 "101000010110101111011100",
						 "101000010110110001101101",
						 "101000010110110011111110",
						 "101000010110110110001111",
						 "101000010110111000100000",
						 "101000010110111010110001",
						 "101000010110111101000010",
						 "101000010110111111010011",
						 "101000010111000001100100",
						 "101000010111000011110101",
						 "101000010111000110000110",
						 "101000010111001000010111",
						 "101000010111001010101000",
						 "101000010111001100111001",
						 "101000010111001111001010",
						 "101000010111010001011011",
						 "101000010110101111011100",
						 "101000010110110001101101",
						 "101000010110110011111110",
						 "101000010110110110001111",
						 "101000010110111000100000",
						 "101000010110111010110001",
						 "101000010110111101000010",
						 "101000010110111111010011",
						 "101000010111000001100100",
						 "101000010111000011110101",
						 "101000010111000110000110",
						 "101000010111001000010111",
						 "101000010111001010101000",
						 "101000010111001100111001",
						 "101000010111001111001010",
						 "101000010111010001011011",
						 "101000010110101111011100",
						 "101000010110110001101100",
						 "101000010110110011111100",
						 "101000010110110110001100",
						 "101000010110111000011100",
						 "101000010110111010101100",
						 "101000010110111100111100",
						 "101000010110111111001100",
						 "101000010111000001011100",
						 "101000010111000011101100",
						 "101000010111000101111100",
						 "101000010111001000001100",
						 "101000010111001010011100",
						 "101000010111001100101100",
						 "101000010111001110111100",
						 "101000010111010001001100",
						 "101000010110101111011100",
						 "101000010110110001101100",
						 "101000010110110011111100",
						 "101000010110110110001100",
						 "101000010110111000011100",
						 "101000010110111010101100",
						 "101000010110111100111100",
						 "101000010110111111001100",
						 "101000010111000001011100",
						 "101000010111000011101100",
						 "101000010111000101111100",
						 "101000010111001000001100",
						 "101000010111001010011100",
						 "101000010111001100101100",
						 "101000010111001110111100",
						 "101000010111010001001100",
						 "101000010110101111011100",
						 "101000010110110001101100",
						 "101000010110110011111100",
						 "101000010110110110001100",
						 "101000010110111000011100",
						 "101000010110111010101100",
						 "101000010110111100111100",
						 "101000010110111111001100",
						 "101000010111000001011100",
						 "101000010111000011101100",
						 "101000010111000101111100",
						 "101000010111001000001100",
						 "101000010111001010011100",
						 "101000010111001100101100",
						 "101000010111001110111100",
						 "101000010111010001001100",
						 "101000011001010010011010",
						 "101000011001010100101001",
						 "101000011001010110111000",
						 "101000011001011001000111",
						 "101000011001011011010110",
						 "101000011001011101100101",
						 "101000011001011111110100",
						 "101000011001100010000011",
						 "101000011001100100010010",
						 "101000011001100110100001",
						 "101000011001101000110000",
						 "101000011001101010111111",
						 "101000011001101101001110",
						 "101000011001101111011101",
						 "101000011001110001101100",
						 "101000011001110011111011",
						 "101000011001010010011010",
						 "101000011001010100101001",
						 "101000011001010110111000",
						 "101000011001011001000111",
						 "101000011001011011010110",
						 "101000011001011101100101",
						 "101000011001011111110100",
						 "101000011001100010000011",
						 "101000011001100100010010",
						 "101000011001100110100001",
						 "101000011001101000110000",
						 "101000011001101010111111",
						 "101000011001101101001110",
						 "101000011001101111011101",
						 "101000011001110001101100",
						 "101000011001110011111011",
						 "101000011001010010011010",
						 "101000011001010100101001",
						 "101000011001010110111000",
						 "101000011001011001000111",
						 "101000011001011011010110",
						 "101000011001011101100101",
						 "101000011001011111110100",
						 "101000011001100010000011",
						 "101000011001100100010010",
						 "101000011001100110100001",
						 "101000011001101000110000",
						 "101000011001101010111111",
						 "101000011001101101001110",
						 "101000011001101111011101",
						 "101000011001110001101100",
						 "101000011001110011111011",
						 "101000011001010010011010",
						 "101000011001010100101000",
						 "101000011001010110110110",
						 "101000011001011001000100",
						 "101000011001011011010010",
						 "101000011001011101100000",
						 "101000011001011111101110",
						 "101000011001100001111100",
						 "101000011001100100001010",
						 "101000011001100110011000",
						 "101000011001101000100110",
						 "101000011001101010110100",
						 "101000011001101101000010",
						 "101000011001101111010000",
						 "101000011001110001011110",
						 "101000011001110011101100",
						 "101000011011110101011000",
						 "101000011011110111100110",
						 "101000011011111001110100",
						 "101000011011111100000010",
						 "101000011011111110010000",
						 "101000011100000000011110",
						 "101000011100000010101100",
						 "101000011100000100111010",
						 "101000011100000111001000",
						 "101000011100001001010110",
						 "101000011100001011100100",
						 "101000011100001101110010",
						 "101000011100010000000000",
						 "101000011100010010001110",
						 "101000011100010100011100",
						 "101000011100010110101010",
						 "101000011011110101011000",
						 "101000011011110111100110",
						 "101000011011111001110100",
						 "101000011011111100000010",
						 "101000011011111110010000",
						 "101000011100000000011110",
						 "101000011100000010101100",
						 "101000011100000100111010",
						 "101000011100000111001000",
						 "101000011100001001010110",
						 "101000011100001011100100",
						 "101000011100001101110010",
						 "101000011100010000000000",
						 "101000011100010010001110",
						 "101000011100010100011100",
						 "101000011100010110101010",
						 "101000011011110101011000",
						 "101000011011110111100110",
						 "101000011011111001110100",
						 "101000011011111100000010",
						 "101000011011111110010000",
						 "101000011100000000011110",
						 "101000011100000010101100",
						 "101000011100000100111010",
						 "101000011100000111001000",
						 "101000011100001001010110",
						 "101000011100001011100100",
						 "101000011100001101110010",
						 "101000011100010000000000",
						 "101000011100010010001110",
						 "101000011100010100011100",
						 "101000011100010110101010",
						 "101000011011110101011000",
						 "101000011011110111100101",
						 "101000011011111001110010",
						 "101000011011111011111111",
						 "101000011011111110001100",
						 "101000011100000000011001",
						 "101000011100000010100110",
						 "101000011100000100110011",
						 "101000011100000111000000",
						 "101000011100001001001101",
						 "101000011100001011011010",
						 "101000011100001101100111",
						 "101000011100001111110100",
						 "101000011100010010000001",
						 "101000011100010100001110",
						 "101000011100010110011011",
						 "101000011011110101011000",
						 "101000011011110111100101",
						 "101000011011111001110010",
						 "101000011011111011111111",
						 "101000011011111110001100",
						 "101000011100000000011001",
						 "101000011100000010100110",
						 "101000011100000100110011",
						 "101000011100000111000000",
						 "101000011100001001001101",
						 "101000011100001011011010",
						 "101000011100001101100111",
						 "101000011100001111110100",
						 "101000011100010010000001",
						 "101000011100010100001110",
						 "101000011100010110011011",
						 "101000011110011000010110",
						 "101000011110011010100011",
						 "101000011110011100110000",
						 "101000011110011110111101",
						 "101000011110100001001010",
						 "101000011110100011010111",
						 "101000011110100101100100",
						 "101000011110100111110001",
						 "101000011110101001111110",
						 "101000011110101100001011",
						 "101000011110101110011000",
						 "101000011110110000100101",
						 "101000011110110010110010",
						 "101000011110110100111111",
						 "101000011110110111001100",
						 "101000011110111001011001",
						 "101000011110011000010110",
						 "101000011110011010100010",
						 "101000011110011100101110",
						 "101000011110011110111010",
						 "101000011110100001000110",
						 "101000011110100011010010",
						 "101000011110100101011110",
						 "101000011110100111101010",
						 "101000011110101001110110",
						 "101000011110101100000010",
						 "101000011110101110001110",
						 "101000011110110000011010",
						 "101000011110110010100110",
						 "101000011110110100110010",
						 "101000011110110110111110",
						 "101000011110111001001010",
						 "101000011110011000010110",
						 "101000011110011010100010",
						 "101000011110011100101110",
						 "101000011110011110111010",
						 "101000011110100001000110",
						 "101000011110100011010010",
						 "101000011110100101011110",
						 "101000011110100111101010",
						 "101000011110101001110110",
						 "101000011110101100000010",
						 "101000011110101110001110",
						 "101000011110110000011010",
						 "101000011110110010100110",
						 "101000011110110100110010",
						 "101000011110110110111110",
						 "101000011110111001001010",
						 "101000011110011000010110",
						 "101000011110011010100010",
						 "101000011110011100101110",
						 "101000011110011110111010",
						 "101000011110100001000110",
						 "101000011110100011010010",
						 "101000011110100101011110",
						 "101000011110100111101010",
						 "101000011110101001110110",
						 "101000011110101100000010",
						 "101000011110101110001110",
						 "101000011110110000011010",
						 "101000011110110010100110",
						 "101000011110110100110010",
						 "101000011110110110111110",
						 "101000011110111001001010",
						 "101000100000111011010100",
						 "101000100000111101011111",
						 "101000100000111111101010",
						 "101000100001000001110101",
						 "101000100001000100000000",
						 "101000100001000110001011",
						 "101000100001001000010110",
						 "101000100001001010100001",
						 "101000100001001100101100",
						 "101000100001001110110111",
						 "101000100001010001000010",
						 "101000100001010011001101",
						 "101000100001010101011000",
						 "101000100001010111100011",
						 "101000100001011001101110",
						 "101000100001011011111001",
						 "101000100000111011010100",
						 "101000100000111101011111",
						 "101000100000111111101010",
						 "101000100001000001110101",
						 "101000100001000100000000",
						 "101000100001000110001011",
						 "101000100001001000010110",
						 "101000100001001010100001",
						 "101000100001001100101100",
						 "101000100001001110110111",
						 "101000100001010001000010",
						 "101000100001010011001101",
						 "101000100001010101011000",
						 "101000100001010111100011",
						 "101000100001011001101110",
						 "101000100001011011111001",
						 "101000100000111011010100",
						 "101000100000111101011111",
						 "101000100000111111101010",
						 "101000100001000001110101",
						 "101000100001000100000000",
						 "101000100001000110001011",
						 "101000100001001000010110",
						 "101000100001001010100001",
						 "101000100001001100101100",
						 "101000100001001110110111",
						 "101000100001010001000010",
						 "101000100001010011001101",
						 "101000100001010101011000",
						 "101000100001010111100011",
						 "101000100001011001101110",
						 "101000100001011011111001",
						 "101000100000111011010100",
						 "101000100000111101011110",
						 "101000100000111111101000",
						 "101000100001000001110010",
						 "101000100001000011111100",
						 "101000100001000110000110",
						 "101000100001001000010000",
						 "101000100001001010011010",
						 "101000100001001100100100",
						 "101000100001001110101110",
						 "101000100001010000111000",
						 "101000100001010011000010",
						 "101000100001010101001100",
						 "101000100001010111010110",
						 "101000100001011001100000",
						 "101000100001011011101010",
						 "101000100000111011010100",
						 "101000100000111101011110",
						 "101000100000111111101000",
						 "101000100001000001110010",
						 "101000100001000011111100",
						 "101000100001000110000110",
						 "101000100001001000010000",
						 "101000100001001010011010",
						 "101000100001001100100100",
						 "101000100001001110101110",
						 "101000100001010000111000",
						 "101000100001010011000010",
						 "101000100001010101001100",
						 "101000100001010111010110",
						 "101000100001011001100000",
						 "101000100001011011101010",
						 "101000100011011110010010",
						 "101000100011100000011100",
						 "101000100011100010100110",
						 "101000100011100100110000",
						 "101000100011100110111010",
						 "101000100011101001000100",
						 "101000100011101011001110",
						 "101000100011101101011000",
						 "101000100011101111100010",
						 "101000100011110001101100",
						 "101000100011110011110110",
						 "101000100011110110000000",
						 "101000100011111000001010",
						 "101000100011111010010100",
						 "101000100011111100011110",
						 "101000100011111110101000",
						 "101000100011011110010010",
						 "101000100011100000011011",
						 "101000100011100010100100",
						 "101000100011100100101101",
						 "101000100011100110110110",
						 "101000100011101000111111",
						 "101000100011101011001000",
						 "101000100011101101010001",
						 "101000100011101111011010",
						 "101000100011110001100011",
						 "101000100011110011101100",
						 "101000100011110101110101",
						 "101000100011110111111110",
						 "101000100011111010000111",
						 "101000100011111100010000",
						 "101000100011111110011001",
						 "101000100011011110010010",
						 "101000100011100000011011",
						 "101000100011100010100100",
						 "101000100011100100101101",
						 "101000100011100110110110",
						 "101000100011101000111111",
						 "101000100011101011001000",
						 "101000100011101101010001",
						 "101000100011101111011010",
						 "101000100011110001100011",
						 "101000100011110011101100",
						 "101000100011110101110101",
						 "101000100011110111111110",
						 "101000100011111010000111",
						 "101000100011111100010000",
						 "101000100011111110011001",
						 "101000100011011110010010",
						 "101000100011100000011011",
						 "101000100011100010100100",
						 "101000100011100100101101",
						 "101000100011100110110110",
						 "101000100011101000111111",
						 "101000100011101011001000",
						 "101000100011101101010001",
						 "101000100011101111011010",
						 "101000100011110001100011",
						 "101000100011110011101100",
						 "101000100011110101110101",
						 "101000100011110111111110",
						 "101000100011111010000111",
						 "101000100011111100010000",
						 "101000100011111110011001",
						 "101000100011011110010010",
						 "101000100011100000011010",
						 "101000100011100010100010",
						 "101000100011100100101010",
						 "101000100011100110110010",
						 "101000100011101000111010",
						 "101000100011101011000010",
						 "101000100011101101001010",
						 "101000100011101111010010",
						 "101000100011110001011010",
						 "101000100011110011100010",
						 "101000100011110101101010",
						 "101000100011110111110010",
						 "101000100011111001111010",
						 "101000100011111100000010",
						 "101000100011111110001010",
						 "101000100110000001010000",
						 "101000100110000011011000",
						 "101000100110000101100000",
						 "101000100110000111101000",
						 "101000100110001001110000",
						 "101000100110001011111000",
						 "101000100110001110000000",
						 "101000100110010000001000",
						 "101000100110010010010000",
						 "101000100110010100011000",
						 "101000100110010110100000",
						 "101000100110011000101000",
						 "101000100110011010110000",
						 "101000100110011100111000",
						 "101000100110011111000000",
						 "101000100110100001001000",
						 "101000100110000001010000",
						 "101000100110000011011000",
						 "101000100110000101100000",
						 "101000100110000111101000",
						 "101000100110001001110000",
						 "101000100110001011111000",
						 "101000100110001110000000",
						 "101000100110010000001000",
						 "101000100110010010010000",
						 "101000100110010100011000",
						 "101000100110010110100000",
						 "101000100110011000101000",
						 "101000100110011010110000",
						 "101000100110011100111000",
						 "101000100110011111000000",
						 "101000100110100001001000",
						 "101000100110000001010000",
						 "101000100110000011010111",
						 "101000100110000101011110",
						 "101000100110000111100101",
						 "101000100110001001101100",
						 "101000100110001011110011",
						 "101000100110001101111010",
						 "101000100110010000000001",
						 "101000100110010010001000",
						 "101000100110010100001111",
						 "101000100110010110010110",
						 "101000100110011000011101",
						 "101000100110011010100100",
						 "101000100110011100101011",
						 "101000100110011110110010",
						 "101000100110100000111001",
						 "101000100110000001010000",
						 "101000100110000011010111",
						 "101000100110000101011110",
						 "101000100110000111100101",
						 "101000100110001001101100",
						 "101000100110001011110011",
						 "101000100110001101111010",
						 "101000100110010000000001",
						 "101000100110010010001000",
						 "101000100110010100001111",
						 "101000100110010110010110",
						 "101000100110011000011101",
						 "101000100110011010100100",
						 "101000100110011100101011",
						 "101000100110011110110010",
						 "101000100110100000111001",
						 "101000100110000001010000",
						 "101000100110000011010111",
						 "101000100110000101011110",
						 "101000100110000111100101",
						 "101000100110001001101100",
						 "101000100110001011110011",
						 "101000100110001101111010",
						 "101000100110010000000001",
						 "101000100110010010001000",
						 "101000100110010100001111",
						 "101000100110010110010110",
						 "101000100110011000011101",
						 "101000100110011010100100",
						 "101000100110011100101011",
						 "101000100110011110110010",
						 "101000100110100000111001",
						 "101000101000100100001110",
						 "101000101000100110010100",
						 "101000101000101000011010",
						 "101000101000101010100000",
						 "101000101000101100100110",
						 "101000101000101110101100",
						 "101000101000110000110010",
						 "101000101000110010111000",
						 "101000101000110100111110",
						 "101000101000110111000100",
						 "101000101000111001001010",
						 "101000101000111011010000",
						 "101000101000111101010110",
						 "101000101000111111011100",
						 "101000101001000001100010",
						 "101000101001000011101000",
						 "101000101000100100001110",
						 "101000101000100110010100",
						 "101000101000101000011010",
						 "101000101000101010100000",
						 "101000101000101100100110",
						 "101000101000101110101100",
						 "101000101000110000110010",
						 "101000101000110010111000",
						 "101000101000110100111110",
						 "101000101000110111000100",
						 "101000101000111001001010",
						 "101000101000111011010000",
						 "101000101000111101010110",
						 "101000101000111111011100",
						 "101000101001000001100010",
						 "101000101001000011101000",
						 "101000101000100100001110",
						 "101000101000100110010100",
						 "101000101000101000011010",
						 "101000101000101010100000",
						 "101000101000101100100110",
						 "101000101000101110101100",
						 "101000101000110000110010",
						 "101000101000110010111000",
						 "101000101000110100111110",
						 "101000101000110111000100",
						 "101000101000111001001010",
						 "101000101000111011010000",
						 "101000101000111101010110",
						 "101000101000111111011100",
						 "101000101001000001100010",
						 "101000101001000011101000",
						 "101000101000100100001110",
						 "101000101000100110010011",
						 "101000101000101000011000",
						 "101000101000101010011101",
						 "101000101000101100100010",
						 "101000101000101110100111",
						 "101000101000110000101100",
						 "101000101000110010110001",
						 "101000101000110100110110",
						 "101000101000110110111011",
						 "101000101000111001000000",
						 "101000101000111011000101",
						 "101000101000111101001010",
						 "101000101000111111001111",
						 "101000101001000001010100",
						 "101000101001000011011001",
						 "101000101011000111001100",
						 "101000101011001001010001",
						 "101000101011001011010110",
						 "101000101011001101011011",
						 "101000101011001111100000",
						 "101000101011010001100101",
						 "101000101011010011101010",
						 "101000101011010101101111",
						 "101000101011010111110100",
						 "101000101011011001111001",
						 "101000101011011011111110",
						 "101000101011011110000011",
						 "101000101011100000001000",
						 "101000101011100010001101",
						 "101000101011100100010010",
						 "101000101011100110010111",
						 "101000101011000111001100",
						 "101000101011001001010001",
						 "101000101011001011010110",
						 "101000101011001101011011",
						 "101000101011001111100000",
						 "101000101011010001100101",
						 "101000101011010011101010",
						 "101000101011010101101111",
						 "101000101011010111110100",
						 "101000101011011001111001",
						 "101000101011011011111110",
						 "101000101011011110000011",
						 "101000101011100000001000",
						 "101000101011100010001101",
						 "101000101011100100010010",
						 "101000101011100110010111",
						 "101000101011000111001100",
						 "101000101011001001010000",
						 "101000101011001011010100",
						 "101000101011001101011000",
						 "101000101011001111011100",
						 "101000101011010001100000",
						 "101000101011010011100100",
						 "101000101011010101101000",
						 "101000101011010111101100",
						 "101000101011011001110000",
						 "101000101011011011110100",
						 "101000101011011101111000",
						 "101000101011011111111100",
						 "101000101011100010000000",
						 "101000101011100100000100",
						 "101000101011100110001000",
						 "101000101011000111001100",
						 "101000101011001001010000",
						 "101000101011001011010100",
						 "101000101011001101011000",
						 "101000101011001111011100",
						 "101000101011010001100000",
						 "101000101011010011100100",
						 "101000101011010101101000",
						 "101000101011010111101100",
						 "101000101011011001110000",
						 "101000101011011011110100",
						 "101000101011011101111000",
						 "101000101011011111111100",
						 "101000101011100010000000",
						 "101000101011100100000100",
						 "101000101011100110001000",
						 "101000101011000111001100",
						 "101000101011001001010000",
						 "101000101011001011010100",
						 "101000101011001101011000",
						 "101000101011001111011100",
						 "101000101011010001100000",
						 "101000101011010011100100",
						 "101000101011010101101000",
						 "101000101011010111101100",
						 "101000101011011001110000",
						 "101000101011011011110100",
						 "101000101011011101111000",
						 "101000101011011111111100",
						 "101000101011100010000000",
						 "101000101011100100000100",
						 "101000101011100110001000",
						 "101000101101101010001010",
						 "101000101101101100001101",
						 "101000101101101110010000",
						 "101000101101110000010011",
						 "101000101101110010010110",
						 "101000101101110100011001",
						 "101000101101110110011100",
						 "101000101101111000011111",
						 "101000101101111010100010",
						 "101000101101111100100101",
						 "101000101101111110101000",
						 "101000101110000000101011",
						 "101000101110000010101110",
						 "101000101110000100110001",
						 "101000101110000110110100",
						 "101000101110001000110111",
						 "101000101101101010001010",
						 "101000101101101100001101",
						 "101000101101101110010000",
						 "101000101101110000010011",
						 "101000101101110010010110",
						 "101000101101110100011001",
						 "101000101101110110011100",
						 "101000101101111000011111",
						 "101000101101111010100010",
						 "101000101101111100100101",
						 "101000101101111110101000",
						 "101000101110000000101011",
						 "101000101110000010101110",
						 "101000101110000100110001",
						 "101000101110000110110100",
						 "101000101110001000110111",
						 "101000101101101010001010",
						 "101000101101101100001101",
						 "101000101101101110010000",
						 "101000101101110000010011",
						 "101000101101110010010110",
						 "101000101101110100011001",
						 "101000101101110110011100",
						 "101000101101111000011111",
						 "101000101101111010100010",
						 "101000101101111100100101",
						 "101000101101111110101000",
						 "101000101110000000101011",
						 "101000101110000010101110",
						 "101000101110000100110001",
						 "101000101110000110110100",
						 "101000101110001000110111",
						 "101000101101101010001010",
						 "101000101101101100001100",
						 "101000101101101110001110",
						 "101000101101110000010000",
						 "101000101101110010010010",
						 "101000101101110100010100",
						 "101000101101110110010110",
						 "101000101101111000011000",
						 "101000101101111010011010",
						 "101000101101111100011100",
						 "101000101101111110011110",
						 "101000101110000000100000",
						 "101000101110000010100010",
						 "101000101110000100100100",
						 "101000101110000110100110",
						 "101000101110001000101000",
						 "101000101101101010001010",
						 "101000101101101100001100",
						 "101000101101101110001110",
						 "101000101101110000010000",
						 "101000101101110010010010",
						 "101000101101110100010100",
						 "101000101101110110010110",
						 "101000101101111000011000",
						 "101000101101111010011010",
						 "101000101101111100011100",
						 "101000101101111110011110",
						 "101000101110000000100000",
						 "101000101110000010100010",
						 "101000101110000100100100",
						 "101000101110000110100110",
						 "101000101110001000101000",
						 "101000110000001101001000",
						 "101000110000001111001010",
						 "101000110000010001001100",
						 "101000110000010011001110",
						 "101000110000010101010000",
						 "101000110000010111010010",
						 "101000110000011001010100",
						 "101000110000011011010110",
						 "101000110000011101011000",
						 "101000110000011111011010",
						 "101000110000100001011100",
						 "101000110000100011011110",
						 "101000110000100101100000",
						 "101000110000100111100010",
						 "101000110000101001100100",
						 "101000110000101011100110",
						 "101000110000001101001000",
						 "101000110000001111001001",
						 "101000110000010001001010",
						 "101000110000010011001011",
						 "101000110000010101001100",
						 "101000110000010111001101",
						 "101000110000011001001110",
						 "101000110000011011001111",
						 "101000110000011101010000",
						 "101000110000011111010001",
						 "101000110000100001010010",
						 "101000110000100011010011",
						 "101000110000100101010100",
						 "101000110000100111010101",
						 "101000110000101001010110",
						 "101000110000101011010111",
						 "101000110000001101001000",
						 "101000110000001111001001",
						 "101000110000010001001010",
						 "101000110000010011001011",
						 "101000110000010101001100",
						 "101000110000010111001101",
						 "101000110000011001001110",
						 "101000110000011011001111",
						 "101000110000011101010000",
						 "101000110000011111010001",
						 "101000110000100001010010",
						 "101000110000100011010011",
						 "101000110000100101010100",
						 "101000110000100111010101",
						 "101000110000101001010110",
						 "101000110000101011010111",
						 "101000110000001101001000",
						 "101000110000001111001001",
						 "101000110000010001001010",
						 "101000110000010011001011",
						 "101000110000010101001100",
						 "101000110000010111001101",
						 "101000110000011001001110",
						 "101000110000011011001111",
						 "101000110000011101010000",
						 "101000110000011111010001",
						 "101000110000100001010010",
						 "101000110000100011010011",
						 "101000110000100101010100",
						 "101000110000100111010101",
						 "101000110000101001010110",
						 "101000110000101011010111",
						 "101000110000001101001000",
						 "101000110000001111001000",
						 "101000110000010001001000",
						 "101000110000010011001000",
						 "101000110000010101001000",
						 "101000110000010111001000",
						 "101000110000011001001000",
						 "101000110000011011001000",
						 "101000110000011101001000",
						 "101000110000011111001000",
						 "101000110000100001001000",
						 "101000110000100011001000",
						 "101000110000100101001000",
						 "101000110000100111001000",
						 "101000110000101001001000",
						 "101000110000101011001000",
						 "101000110010110000000110",
						 "101000110010110010000110",
						 "101000110010110100000110",
						 "101000110010110110000110",
						 "101000110010111000000110",
						 "101000110010111010000110",
						 "101000110010111100000110",
						 "101000110010111110000110",
						 "101000110011000000000110",
						 "101000110011000010000110",
						 "101000110011000100000110",
						 "101000110011000110000110",
						 "101000110011001000000110",
						 "101000110011001010000110",
						 "101000110011001100000110",
						 "101000110011001110000110",
						 "101000110010110000000110",
						 "101000110010110010000110",
						 "101000110010110100000110",
						 "101000110010110110000110",
						 "101000110010111000000110",
						 "101000110010111010000110",
						 "101000110010111100000110",
						 "101000110010111110000110",
						 "101000110011000000000110",
						 "101000110011000010000110",
						 "101000110011000100000110",
						 "101000110011000110000110",
						 "101000110011001000000110",
						 "101000110011001010000110",
						 "101000110011001100000110",
						 "101000110011001110000110",
						 "101000110010110000000110",
						 "101000110010110010000101",
						 "101000110010110100000100",
						 "101000110010110110000011",
						 "101000110010111000000010",
						 "101000110010111010000001",
						 "101000110010111100000000",
						 "101000110010111101111111",
						 "101000110010111111111110",
						 "101000110011000001111101",
						 "101000110011000011111100",
						 "101000110011000101111011",
						 "101000110011000111111010",
						 "101000110011001001111001",
						 "101000110011001011111000",
						 "101000110011001101110111",
						 "101000110010110000000110",
						 "101000110010110010000101",
						 "101000110010110100000100",
						 "101000110010110110000011",
						 "101000110010111000000010",
						 "101000110010111010000001",
						 "101000110010111100000000",
						 "101000110010111101111111",
						 "101000110010111111111110",
						 "101000110011000001111101",
						 "101000110011000011111100",
						 "101000110011000101111011",
						 "101000110011000111111010",
						 "101000110011001001111001",
						 "101000110011001011111000",
						 "101000110011001101110111",
						 "101000110010110000000110",
						 "101000110010110010000101",
						 "101000110010110100000100",
						 "101000110010110110000011",
						 "101000110010111000000010",
						 "101000110010111010000001",
						 "101000110010111100000000",
						 "101000110010111101111111",
						 "101000110010111111111110",
						 "101000110011000001111101",
						 "101000110011000011111100",
						 "101000110011000101111011",
						 "101000110011000111111010",
						 "101000110011001001111001",
						 "101000110011001011111000",
						 "101000110011001101110111",
						 "101000110010110000000110",
						 "101000110010110010000100",
						 "101000110010110100000010",
						 "101000110010110110000000",
						 "101000110010110111111110",
						 "101000110010111001111100",
						 "101000110010111011111010",
						 "101000110010111101111000",
						 "101000110010111111110110",
						 "101000110011000001110100",
						 "101000110011000011110010",
						 "101000110011000101110000",
						 "101000110011000111101110",
						 "101000110011001001101100",
						 "101000110011001011101010",
						 "101000110011001101101000",
						 "101000110101010011000100",
						 "101000110101010101000010",
						 "101000110101010111000000",
						 "101000110101011000111110",
						 "101000110101011010111100",
						 "101000110101011100111010",
						 "101000110101011110111000",
						 "101000110101100000110110",
						 "101000110101100010110100",
						 "101000110101100100110010",
						 "101000110101100110110000",
						 "101000110101101000101110",
						 "101000110101101010101100",
						 "101000110101101100101010",
						 "101000110101101110101000",
						 "101000110101110000100110",
						 "101000110101010011000100",
						 "101000110101010101000010",
						 "101000110101010111000000",
						 "101000110101011000111110",
						 "101000110101011010111100",
						 "101000110101011100111010",
						 "101000110101011110111000",
						 "101000110101100000110110",
						 "101000110101100010110100",
						 "101000110101100100110010",
						 "101000110101100110110000",
						 "101000110101101000101110",
						 "101000110101101010101100",
						 "101000110101101100101010",
						 "101000110101101110101000",
						 "101000110101110000100110",
						 "101000110101010011000100",
						 "101000110101010101000001",
						 "101000110101010110111110",
						 "101000110101011000111011",
						 "101000110101011010111000",
						 "101000110101011100110101",
						 "101000110101011110110010",
						 "101000110101100000101111",
						 "101000110101100010101100",
						 "101000110101100100101001",
						 "101000110101100110100110",
						 "101000110101101000100011",
						 "101000110101101010100000",
						 "101000110101101100011101",
						 "101000110101101110011010",
						 "101000110101110000010111",
						 "101000110101010011000100",
						 "101000110101010101000001",
						 "101000110101010110111110",
						 "101000110101011000111011",
						 "101000110101011010111000",
						 "101000110101011100110101",
						 "101000110101011110110010",
						 "101000110101100000101111",
						 "101000110101100010101100",
						 "101000110101100100101001",
						 "101000110101100110100110",
						 "101000110101101000100011",
						 "101000110101101010100000",
						 "101000110101101100011101",
						 "101000110101101110011010",
						 "101000110101110000010111",
						 "101000110101010011000100",
						 "101000110101010101000000",
						 "101000110101010110111100",
						 "101000110101011000111000",
						 "101000110101011010110100",
						 "101000110101011100110000",
						 "101000110101011110101100",
						 "101000110101100000101000",
						 "101000110101100010100100",
						 "101000110101100100100000",
						 "101000110101100110011100",
						 "101000110101101000011000",
						 "101000110101101010010100",
						 "101000110101101100010000",
						 "101000110101101110001100",
						 "101000110101110000001000",
						 "101000110111110110000010",
						 "101000110111110111111110",
						 "101000110111111001111010",
						 "101000110111111011110110",
						 "101000110111111101110010",
						 "101000110111111111101110",
						 "101000111000000001101010",
						 "101000111000000011100110",
						 "101000111000000101100010",
						 "101000111000000111011110",
						 "101000111000001001011010",
						 "101000111000001011010110",
						 "101000111000001101010010",
						 "101000111000001111001110",
						 "101000111000010001001010",
						 "101000111000010011000110",
						 "101000110111110110000010",
						 "101000110111110111111110",
						 "101000110111111001111010",
						 "101000110111111011110110",
						 "101000110111111101110010",
						 "101000110111111111101110",
						 "101000111000000001101010",
						 "101000111000000011100110",
						 "101000111000000101100010",
						 "101000111000000111011110",
						 "101000111000001001011010",
						 "101000111000001011010110",
						 "101000111000001101010010",
						 "101000111000001111001110",
						 "101000111000010001001010",
						 "101000111000010011000110",
						 "101000110111110110000010",
						 "101000110111110111111101",
						 "101000110111111001111000",
						 "101000110111111011110011",
						 "101000110111111101101110",
						 "101000110111111111101001",
						 "101000111000000001100100",
						 "101000111000000011011111",
						 "101000111000000101011010",
						 "101000111000000111010101",
						 "101000111000001001010000",
						 "101000111000001011001011",
						 "101000111000001101000110",
						 "101000111000001111000001",
						 "101000111000010000111100",
						 "101000111000010010110111",
						 "101000110111110110000010",
						 "101000110111110111111101",
						 "101000110111111001111000",
						 "101000110111111011110011",
						 "101000110111111101101110",
						 "101000110111111111101001",
						 "101000111000000001100100",
						 "101000111000000011011111",
						 "101000111000000101011010",
						 "101000111000000111010101",
						 "101000111000001001010000",
						 "101000111000001011001011",
						 "101000111000001101000110",
						 "101000111000001111000001",
						 "101000111000010000111100",
						 "101000111000010010110111",
						 "101000110111110110000010",
						 "101000110111110111111101",
						 "101000110111111001111000",
						 "101000110111111011110011",
						 "101000110111111101101110",
						 "101000110111111111101001",
						 "101000111000000001100100",
						 "101000111000000011011111",
						 "101000111000000101011010",
						 "101000111000000111010101",
						 "101000111000001001010000",
						 "101000111000001011001011",
						 "101000111000001101000110",
						 "101000111000001111000001",
						 "101000111000010000111100",
						 "101000111000010010110111",
						 "101000111010011001000000",
						 "101000111010011010111010",
						 "101000111010011100110100",
						 "101000111010011110101110",
						 "101000111010100000101000",
						 "101000111010100010100010",
						 "101000111010100100011100",
						 "101000111010100110010110",
						 "101000111010101000010000",
						 "101000111010101010001010",
						 "101000111010101100000100",
						 "101000111010101101111110",
						 "101000111010101111111000",
						 "101000111010110001110010",
						 "101000111010110011101100",
						 "101000111010110101100110",
						 "101000111010011001000000",
						 "101000111010011010111010",
						 "101000111010011100110100",
						 "101000111010011110101110",
						 "101000111010100000101000",
						 "101000111010100010100010",
						 "101000111010100100011100",
						 "101000111010100110010110",
						 "101000111010101000010000",
						 "101000111010101010001010",
						 "101000111010101100000100",
						 "101000111010101101111110",
						 "101000111010101111111000",
						 "101000111010110001110010",
						 "101000111010110011101100",
						 "101000111010110101100110",
						 "101000111010011001000000",
						 "101000111010011010111010",
						 "101000111010011100110100",
						 "101000111010011110101110",
						 "101000111010100000101000",
						 "101000111010100010100010",
						 "101000111010100100011100",
						 "101000111010100110010110",
						 "101000111010101000010000",
						 "101000111010101010001010",
						 "101000111010101100000100",
						 "101000111010101101111110",
						 "101000111010101111111000",
						 "101000111010110001110010",
						 "101000111010110011101100",
						 "101000111010110101100110",
						 "101000111010011001000000",
						 "101000111010011010111001",
						 "101000111010011100110010",
						 "101000111010011110101011",
						 "101000111010100000100100",
						 "101000111010100010011101",
						 "101000111010100100010110",
						 "101000111010100110001111",
						 "101000111010101000001000",
						 "101000111010101010000001",
						 "101000111010101011111010",
						 "101000111010101101110011",
						 "101000111010101111101100",
						 "101000111010110001100101",
						 "101000111010110011011110",
						 "101000111010110101010111",
						 "101000111010011001000000",
						 "101000111010011010111001",
						 "101000111010011100110010",
						 "101000111010011110101011",
						 "101000111010100000100100",
						 "101000111010100010011101",
						 "101000111010100100010110",
						 "101000111010100110001111",
						 "101000111010101000001000",
						 "101000111010101010000001",
						 "101000111010101011111010",
						 "101000111010101101110011",
						 "101000111010101111101100",
						 "101000111010110001100101",
						 "101000111010110011011110",
						 "101000111010110101010111",
						 "101000111100111011111110",
						 "101000111100111101110111",
						 "101000111100111111110000",
						 "101000111101000001101001",
						 "101000111101000011100010",
						 "101000111101000101011011",
						 "101000111101000111010100",
						 "101000111101001001001101",
						 "101000111101001011000110",
						 "101000111101001100111111",
						 "101000111101001110111000",
						 "101000111101010000110001",
						 "101000111101010010101010",
						 "101000111101010100100011",
						 "101000111101010110011100",
						 "101000111101011000010101",
						 "101000111100111011111110",
						 "101000111100111101110110",
						 "101000111100111111101110",
						 "101000111101000001100110",
						 "101000111101000011011110",
						 "101000111101000101010110",
						 "101000111101000111001110",
						 "101000111101001001000110",
						 "101000111101001010111110",
						 "101000111101001100110110",
						 "101000111101001110101110",
						 "101000111101010000100110",
						 "101000111101010010011110",
						 "101000111101010100010110",
						 "101000111101010110001110",
						 "101000111101011000000110",
						 "101000111100111011111110",
						 "101000111100111101110110",
						 "101000111100111111101110",
						 "101000111101000001100110",
						 "101000111101000011011110",
						 "101000111101000101010110",
						 "101000111101000111001110",
						 "101000111101001001000110",
						 "101000111101001010111110",
						 "101000111101001100110110",
						 "101000111101001110101110",
						 "101000111101010000100110",
						 "101000111101010010011110",
						 "101000111101010100010110",
						 "101000111101010110001110",
						 "101000111101011000000110",
						 "101000111100111011111110",
						 "101000111100111101110110",
						 "101000111100111111101110",
						 "101000111101000001100110",
						 "101000111101000011011110",
						 "101000111101000101010110",
						 "101000111101000111001110",
						 "101000111101001001000110",
						 "101000111101001010111110",
						 "101000111101001100110110",
						 "101000111101001110101110",
						 "101000111101010000100110",
						 "101000111101010010011110",
						 "101000111101010100010110",
						 "101000111101010110001110",
						 "101000111101011000000110",
						 "101000111100111011111110",
						 "101000111100111101110101",
						 "101000111100111111101100",
						 "101000111101000001100011",
						 "101000111101000011011010",
						 "101000111101000101010001",
						 "101000111101000111001000",
						 "101000111101001000111111",
						 "101000111101001010110110",
						 "101000111101001100101101",
						 "101000111101001110100100",
						 "101000111101010000011011",
						 "101000111101010010010010",
						 "101000111101010100001001",
						 "101000111101010110000000",
						 "101000111101010111110111",
						 "101000111100111011111110",
						 "101000111100111101110101",
						 "101000111100111111101100",
						 "101000111101000001100011",
						 "101000111101000011011010",
						 "101000111101000101010001",
						 "101000111101000111001000",
						 "101000111101001000111111",
						 "101000111101001010110110",
						 "101000111101001100101101",
						 "101000111101001110100100",
						 "101000111101010000011011",
						 "101000111101010010010010",
						 "101000111101010100001001",
						 "101000111101010110000000",
						 "101000111101010111110111",
						 "101000111111011110111100",
						 "101000111111100000110011",
						 "101000111111100010101010",
						 "101000111111100100100001",
						 "101000111111100110011000",
						 "101000111111101000001111",
						 "101000111111101010000110",
						 "101000111111101011111101",
						 "101000111111101101110100",
						 "101000111111101111101011",
						 "101000111111110001100010",
						 "101000111111110011011001",
						 "101000111111110101010000",
						 "101000111111110111000111",
						 "101000111111111000111110",
						 "101000111111111010110101",
						 "101000111111011110111100",
						 "101000111111100000110010",
						 "101000111111100010101000",
						 "101000111111100100011110",
						 "101000111111100110010100",
						 "101000111111101000001010",
						 "101000111111101010000000",
						 "101000111111101011110110",
						 "101000111111101101101100",
						 "101000111111101111100010",
						 "101000111111110001011000",
						 "101000111111110011001110",
						 "101000111111110101000100",
						 "101000111111110110111010",
						 "101000111111111000110000",
						 "101000111111111010100110",
						 "101000111111011110111100",
						 "101000111111100000110010",
						 "101000111111100010101000",
						 "101000111111100100011110",
						 "101000111111100110010100",
						 "101000111111101000001010",
						 "101000111111101010000000",
						 "101000111111101011110110",
						 "101000111111101101101100",
						 "101000111111101111100010",
						 "101000111111110001011000",
						 "101000111111110011001110",
						 "101000111111110101000100",
						 "101000111111110110111010",
						 "101000111111111000110000",
						 "101000111111111010100110",
						 "101000111111011110111100",
						 "101000111111100000110010",
						 "101000111111100010101000",
						 "101000111111100100011110",
						 "101000111111100110010100",
						 "101000111111101000001010",
						 "101000111111101010000000",
						 "101000111111101011110110",
						 "101000111111101101101100",
						 "101000111111101111100010",
						 "101000111111110001011000",
						 "101000111111110011001110",
						 "101000111111110101000100",
						 "101000111111110110111010",
						 "101000111111111000110000",
						 "101000111111111010100110",
						 "101000111111011110111100",
						 "101000111111100000110001",
						 "101000111111100010100110",
						 "101000111111100100011011",
						 "101000111111100110010000",
						 "101000111111101000000101",
						 "101000111111101001111010",
						 "101000111111101011101111",
						 "101000111111101101100100",
						 "101000111111101111011001",
						 "101000111111110001001110",
						 "101000111111110011000011",
						 "101000111111110100111000",
						 "101000111111110110101101",
						 "101000111111111000100010",
						 "101000111111111010010111",
						 "101001000010000001111010",
						 "101001000010000011101111",
						 "101001000010000101100100",
						 "101001000010000111011001",
						 "101001000010001001001110",
						 "101001000010001011000011",
						 "101001000010001100111000",
						 "101001000010001110101101",
						 "101001000010010000100010",
						 "101001000010010010010111",
						 "101001000010010100001100",
						 "101001000010010110000001",
						 "101001000010010111110110",
						 "101001000010011001101011",
						 "101001000010011011100000",
						 "101001000010011101010101",
						 "101001000010000001111010",
						 "101001000010000011101111",
						 "101001000010000101100100",
						 "101001000010000111011001",
						 "101001000010001001001110",
						 "101001000010001011000011",
						 "101001000010001100111000",
						 "101001000010001110101101",
						 "101001000010010000100010",
						 "101001000010010010010111",
						 "101001000010010100001100",
						 "101001000010010110000001",
						 "101001000010010111110110",
						 "101001000010011001101011",
						 "101001000010011011100000",
						 "101001000010011101010101",
						 "101001000010000001111010",
						 "101001000010000011101110",
						 "101001000010000101100010",
						 "101001000010000111010110",
						 "101001000010001001001010",
						 "101001000010001010111110",
						 "101001000010001100110010",
						 "101001000010001110100110",
						 "101001000010010000011010",
						 "101001000010010010001110",
						 "101001000010010100000010",
						 "101001000010010101110110",
						 "101001000010010111101010",
						 "101001000010011001011110",
						 "101001000010011011010010",
						 "101001000010011101000110",
						 "101001000010000001111010",
						 "101001000010000011101110",
						 "101001000010000101100010",
						 "101001000010000111010110",
						 "101001000010001001001010",
						 "101001000010001010111110",
						 "101001000010001100110010",
						 "101001000010001110100110",
						 "101001000010010000011010",
						 "101001000010010010001110",
						 "101001000010010100000010",
						 "101001000010010101110110",
						 "101001000010010111101010",
						 "101001000010011001011110",
						 "101001000010011011010010",
						 "101001000010011101000110",
						 "101001000010000001111010",
						 "101001000010000011101110",
						 "101001000010000101100010",
						 "101001000010000111010110",
						 "101001000010001001001010",
						 "101001000010001010111110",
						 "101001000010001100110010",
						 "101001000010001110100110",
						 "101001000010010000011010",
						 "101001000010010010001110",
						 "101001000010010100000010",
						 "101001000010010101110110",
						 "101001000010010111101010",
						 "101001000010011001011110",
						 "101001000010011011010010",
						 "101001000010011101000110",
						 "101001000010000001111010",
						 "101001000010000011101101",
						 "101001000010000101100000",
						 "101001000010000111010011",
						 "101001000010001001000110",
						 "101001000010001010111001",
						 "101001000010001100101100",
						 "101001000010001110011111",
						 "101001000010010000010010",
						 "101001000010010010000101",
						 "101001000010010011111000",
						 "101001000010010101101011",
						 "101001000010010111011110",
						 "101001000010011001010001",
						 "101001000010011011000100",
						 "101001000010011100110111",
						 "101001000100100100111000",
						 "101001000100100110101011",
						 "101001000100101000011110",
						 "101001000100101010010001",
						 "101001000100101100000100",
						 "101001000100101101110111",
						 "101001000100101111101010",
						 "101001000100110001011101",
						 "101001000100110011010000",
						 "101001000100110101000011",
						 "101001000100110110110110",
						 "101001000100111000101001",
						 "101001000100111010011100",
						 "101001000100111100001111",
						 "101001000100111110000010",
						 "101001000100111111110101",
						 "101001000100100100111000",
						 "101001000100100110101010",
						 "101001000100101000011100",
						 "101001000100101010001110",
						 "101001000100101100000000",
						 "101001000100101101110010",
						 "101001000100101111100100",
						 "101001000100110001010110",
						 "101001000100110011001000",
						 "101001000100110100111010",
						 "101001000100110110101100",
						 "101001000100111000011110",
						 "101001000100111010010000",
						 "101001000100111100000010",
						 "101001000100111101110100",
						 "101001000100111111100110",
						 "101001000100100100111000",
						 "101001000100100110101010",
						 "101001000100101000011100",
						 "101001000100101010001110",
						 "101001000100101100000000",
						 "101001000100101101110010",
						 "101001000100101111100100",
						 "101001000100110001010110",
						 "101001000100110011001000",
						 "101001000100110100111010",
						 "101001000100110110101100",
						 "101001000100111000011110",
						 "101001000100111010010000",
						 "101001000100111100000010",
						 "101001000100111101110100",
						 "101001000100111111100110",
						 "101001000100100100111000",
						 "101001000100100110101010",
						 "101001000100101000011100",
						 "101001000100101010001110",
						 "101001000100101100000000",
						 "101001000100101101110010",
						 "101001000100101111100100",
						 "101001000100110001010110",
						 "101001000100110011001000",
						 "101001000100110100111010",
						 "101001000100110110101100",
						 "101001000100111000011110",
						 "101001000100111010010000",
						 "101001000100111100000010",
						 "101001000100111101110100",
						 "101001000100111111100110",
						 "101001000100100100111000",
						 "101001000100100110101001",
						 "101001000100101000011010",
						 "101001000100101010001011",
						 "101001000100101011111100",
						 "101001000100101101101101",
						 "101001000100101111011110",
						 "101001000100110001001111",
						 "101001000100110011000000",
						 "101001000100110100110001",
						 "101001000100110110100010",
						 "101001000100111000010011",
						 "101001000100111010000100",
						 "101001000100111011110101",
						 "101001000100111101100110",
						 "101001000100111111010111",
						 "101001000100100100111000",
						 "101001000100100110101001",
						 "101001000100101000011010",
						 "101001000100101010001011",
						 "101001000100101011111100",
						 "101001000100101101101101",
						 "101001000100101111011110",
						 "101001000100110001001111",
						 "101001000100110011000000",
						 "101001000100110100110001",
						 "101001000100110110100010",
						 "101001000100111000010011",
						 "101001000100111010000100",
						 "101001000100111011110101",
						 "101001000100111101100110",
						 "101001000100111111010111",
						 "101001000111000111110110",
						 "101001000111001001100111",
						 "101001000111001011011000",
						 "101001000111001101001001",
						 "101001000111001110111010",
						 "101001000111010000101011",
						 "101001000111010010011100",
						 "101001000111010100001101",
						 "101001000111010101111110",
						 "101001000111010111101111",
						 "101001000111011001100000",
						 "101001000111011011010001",
						 "101001000111011101000010",
						 "101001000111011110110011",
						 "101001000111100000100100",
						 "101001000111100010010101",
						 "101001000111000111110110",
						 "101001000111001001100110",
						 "101001000111001011010110",
						 "101001000111001101000110",
						 "101001000111001110110110",
						 "101001000111010000100110",
						 "101001000111010010010110",
						 "101001000111010100000110",
						 "101001000111010101110110",
						 "101001000111010111100110",
						 "101001000111011001010110",
						 "101001000111011011000110",
						 "101001000111011100110110",
						 "101001000111011110100110",
						 "101001000111100000010110",
						 "101001000111100010000110",
						 "101001000111000111110110",
						 "101001000111001001100110",
						 "101001000111001011010110",
						 "101001000111001101000110",
						 "101001000111001110110110",
						 "101001000111010000100110",
						 "101001000111010010010110",
						 "101001000111010100000110",
						 "101001000111010101110110",
						 "101001000111010111100110",
						 "101001000111011001010110",
						 "101001000111011011000110",
						 "101001000111011100110110",
						 "101001000111011110100110",
						 "101001000111100000010110",
						 "101001000111100010000110",
						 "101001000111000111110110",
						 "101001000111001001100110",
						 "101001000111001011010110",
						 "101001000111001101000110",
						 "101001000111001110110110",
						 "101001000111010000100110",
						 "101001000111010010010110",
						 "101001000111010100000110",
						 "101001000111010101110110",
						 "101001000111010111100110",
						 "101001000111011001010110",
						 "101001000111011011000110",
						 "101001000111011100110110",
						 "101001000111011110100110",
						 "101001000111100000010110",
						 "101001000111100010000110",
						 "101001000111000111110110",
						 "101001000111001001100101",
						 "101001000111001011010100",
						 "101001000111001101000011",
						 "101001000111001110110010",
						 "101001000111010000100001",
						 "101001000111010010010000",
						 "101001000111010011111111",
						 "101001000111010101101110",
						 "101001000111010111011101",
						 "101001000111011001001100",
						 "101001000111011010111011",
						 "101001000111011100101010",
						 "101001000111011110011001",
						 "101001000111100000001000",
						 "101001000111100001110111",
						 "101001001001101010110100",
						 "101001001001101100100011",
						 "101001001001101110010010",
						 "101001001001110000000001",
						 "101001001001110001110000",
						 "101001001001110011011111",
						 "101001001001110101001110",
						 "101001001001110110111101",
						 "101001001001111000101100",
						 "101001001001111010011011",
						 "101001001001111100001010",
						 "101001001001111101111001",
						 "101001001001111111101000",
						 "101001001010000001010111",
						 "101001001010000011000110",
						 "101001001010000100110101",
						 "101001001001101010110100",
						 "101001001001101100100011",
						 "101001001001101110010010",
						 "101001001001110000000001",
						 "101001001001110001110000",
						 "101001001001110011011111",
						 "101001001001110101001110",
						 "101001001001110110111101",
						 "101001001001111000101100",
						 "101001001001111010011011",
						 "101001001001111100001010",
						 "101001001001111101111001",
						 "101001001001111111101000",
						 "101001001010000001010111",
						 "101001001010000011000110",
						 "101001001010000100110101",
						 "101001001001101010110100",
						 "101001001001101100100010",
						 "101001001001101110010000",
						 "101001001001101111111110",
						 "101001001001110001101100",
						 "101001001001110011011010",
						 "101001001001110101001000",
						 "101001001001110110110110",
						 "101001001001111000100100",
						 "101001001001111010010010",
						 "101001001001111100000000",
						 "101001001001111101101110",
						 "101001001001111111011100",
						 "101001001010000001001010",
						 "101001001010000010111000",
						 "101001001010000100100110",
						 "101001001001101010110100",
						 "101001001001101100100010",
						 "101001001001101110010000",
						 "101001001001101111111110",
						 "101001001001110001101100",
						 "101001001001110011011010",
						 "101001001001110101001000",
						 "101001001001110110110110",
						 "101001001001111000100100",
						 "101001001001111010010010",
						 "101001001001111100000000",
						 "101001001001111101101110",
						 "101001001001111111011100",
						 "101001001010000001001010",
						 "101001001010000010111000",
						 "101001001010000100100110",
						 "101001001001101010110100",
						 "101001001001101100100010",
						 "101001001001101110010000",
						 "101001001001101111111110",
						 "101001001001110001101100",
						 "101001001001110011011010",
						 "101001001001110101001000",
						 "101001001001110110110110",
						 "101001001001111000100100",
						 "101001001001111010010010",
						 "101001001001111100000000",
						 "101001001001111101101110",
						 "101001001001111111011100",
						 "101001001010000001001010",
						 "101001001010000010111000",
						 "101001001010000100100110",
						 "101001001001101010110100",
						 "101001001001101100100001",
						 "101001001001101110001110",
						 "101001001001101111111011",
						 "101001001001110001101000",
						 "101001001001110011010101",
						 "101001001001110101000010",
						 "101001001001110110101111",
						 "101001001001111000011100",
						 "101001001001111010001001",
						 "101001001001111011110110",
						 "101001001001111101100011",
						 "101001001001111111010000",
						 "101001001010000000111101",
						 "101001001010000010101010",
						 "101001001010000100010111",
						 "101001001100001101110010",
						 "101001001100001111011111",
						 "101001001100010001001100",
						 "101001001100010010111001",
						 "101001001100010100100110",
						 "101001001100010110010011",
						 "101001001100011000000000",
						 "101001001100011001101101",
						 "101001001100011011011010",
						 "101001001100011101000111",
						 "101001001100011110110100",
						 "101001001100100000100001",
						 "101001001100100010001110",
						 "101001001100100011111011",
						 "101001001100100101101000",
						 "101001001100100111010101",
						 "101001001100001101110010",
						 "101001001100001111011110",
						 "101001001100010001001010",
						 "101001001100010010110110",
						 "101001001100010100100010",
						 "101001001100010110001110",
						 "101001001100010111111010",
						 "101001001100011001100110",
						 "101001001100011011010010",
						 "101001001100011100111110",
						 "101001001100011110101010",
						 "101001001100100000010110",
						 "101001001100100010000010",
						 "101001001100100011101110",
						 "101001001100100101011010",
						 "101001001100100111000110",
						 "101001001100001101110010",
						 "101001001100001111011110",
						 "101001001100010001001010",
						 "101001001100010010110110",
						 "101001001100010100100010",
						 "101001001100010110001110",
						 "101001001100010111111010",
						 "101001001100011001100110",
						 "101001001100011011010010",
						 "101001001100011100111110",
						 "101001001100011110101010",
						 "101001001100100000010110",
						 "101001001100100010000010",
						 "101001001100100011101110",
						 "101001001100100101011010",
						 "101001001100100111000110",
						 "101001001100001101110010",
						 "101001001100001111011110",
						 "101001001100010001001010",
						 "101001001100010010110110",
						 "101001001100010100100010",
						 "101001001100010110001110",
						 "101001001100010111111010",
						 "101001001100011001100110",
						 "101001001100011011010010",
						 "101001001100011100111110",
						 "101001001100011110101010",
						 "101001001100100000010110",
						 "101001001100100010000010",
						 "101001001100100011101110",
						 "101001001100100101011010",
						 "101001001100100111000110",
						 "101001001100001101110010",
						 "101001001100001111011101",
						 "101001001100010001001000",
						 "101001001100010010110011",
						 "101001001100010100011110",
						 "101001001100010110001001",
						 "101001001100010111110100",
						 "101001001100011001011111",
						 "101001001100011011001010",
						 "101001001100011100110101",
						 "101001001100011110100000",
						 "101001001100100000001011",
						 "101001001100100001110110",
						 "101001001100100011100001",
						 "101001001100100101001100",
						 "101001001100100110110111",
						 "101001001100001101110010",
						 "101001001100001111011101",
						 "101001001100010001001000",
						 "101001001100010010110011",
						 "101001001100010100011110",
						 "101001001100010110001001",
						 "101001001100010111110100",
						 "101001001100011001011111",
						 "101001001100011011001010",
						 "101001001100011100110101",
						 "101001001100011110100000",
						 "101001001100100000001011",
						 "101001001100100001110110",
						 "101001001100100011100001",
						 "101001001100100101001100",
						 "101001001100100110110111",
						 "101001001110110000110000",
						 "101001001110110010011011",
						 "101001001110110100000110",
						 "101001001110110101110001",
						 "101001001110110111011100",
						 "101001001110111001000111",
						 "101001001110111010110010",
						 "101001001110111100011101",
						 "101001001110111110001000",
						 "101001001110111111110011",
						 "101001001111000001011110",
						 "101001001111000011001001",
						 "101001001111000100110100",
						 "101001001111000110011111",
						 "101001001111001000001010",
						 "101001001111001001110101",
						 "101001001110110000110000",
						 "101001001110110010011010",
						 "101001001110110100000100",
						 "101001001110110101101110",
						 "101001001110110111011000",
						 "101001001110111001000010",
						 "101001001110111010101100",
						 "101001001110111100010110",
						 "101001001110111110000000",
						 "101001001110111111101010",
						 "101001001111000001010100",
						 "101001001111000010111110",
						 "101001001111000100101000",
						 "101001001111000110010010",
						 "101001001111000111111100",
						 "101001001111001001100110",
						 "101001001110110000110000",
						 "101001001110110010011010",
						 "101001001110110100000100",
						 "101001001110110101101110",
						 "101001001110110111011000",
						 "101001001110111001000010",
						 "101001001110111010101100",
						 "101001001110111100010110",
						 "101001001110111110000000",
						 "101001001110111111101010",
						 "101001001111000001010100",
						 "101001001111000010111110",
						 "101001001111000100101000",
						 "101001001111000110010010",
						 "101001001111000111111100",
						 "101001001111001001100110",
						 "101001001110110000110000",
						 "101001001110110010011010",
						 "101001001110110100000100",
						 "101001001110110101101110",
						 "101001001110110111011000",
						 "101001001110111001000010",
						 "101001001110111010101100",
						 "101001001110111100010110",
						 "101001001110111110000000",
						 "101001001110111111101010",
						 "101001001111000001010100",
						 "101001001111000010111110",
						 "101001001111000100101000",
						 "101001001111000110010010",
						 "101001001111000111111100",
						 "101001001111001001100110",
						 "101001001110110000110000",
						 "101001001110110010011001",
						 "101001001110110100000010",
						 "101001001110110101101011",
						 "101001001110110111010100",
						 "101001001110111000111101",
						 "101001001110111010100110",
						 "101001001110111100001111",
						 "101001001110111101111000",
						 "101001001110111111100001",
						 "101001001111000001001010",
						 "101001001111000010110011",
						 "101001001111000100011100",
						 "101001001111000110000101",
						 "101001001111000111101110",
						 "101001001111001001010111",
						 "101001001110110000110000",
						 "101001001110110010011001",
						 "101001001110110100000010",
						 "101001001110110101101011",
						 "101001001110110111010100",
						 "101001001110111000111101",
						 "101001001110111010100110",
						 "101001001110111100001111",
						 "101001001110111101111000",
						 "101001001110111111100001",
						 "101001001111000001001010",
						 "101001001111000010110011",
						 "101001001111000100011100",
						 "101001001111000110000101",
						 "101001001111000111101110",
						 "101001001111001001010111",
						 "101001001110110000110000",
						 "101001001110110010011001",
						 "101001001110110100000010",
						 "101001001110110101101011",
						 "101001001110110111010100",
						 "101001001110111000111101",
						 "101001001110111010100110",
						 "101001001110111100001111",
						 "101001001110111101111000",
						 "101001001110111111100001",
						 "101001001111000001001010",
						 "101001001111000010110011",
						 "101001001111000100011100",
						 "101001001111000110000101",
						 "101001001111000111101110",
						 "101001001111001001010111",
						 "101001010001010011101110",
						 "101001010001010101010110",
						 "101001010001010110111110",
						 "101001010001011000100110",
						 "101001010001011010001110",
						 "101001010001011011110110",
						 "101001010001011101011110",
						 "101001010001011111000110",
						 "101001010001100000101110",
						 "101001010001100010010110",
						 "101001010001100011111110",
						 "101001010001100101100110",
						 "101001010001100111001110",
						 "101001010001101000110110",
						 "101001010001101010011110",
						 "101001010001101100000110",
						 "101001010001010011101110",
						 "101001010001010101010110",
						 "101001010001010110111110",
						 "101001010001011000100110",
						 "101001010001011010001110",
						 "101001010001011011110110",
						 "101001010001011101011110",
						 "101001010001011111000110",
						 "101001010001100000101110",
						 "101001010001100010010110",
						 "101001010001100011111110",
						 "101001010001100101100110",
						 "101001010001100111001110",
						 "101001010001101000110110",
						 "101001010001101010011110",
						 "101001010001101100000110",
						 "101001010001010011101110",
						 "101001010001010101010110",
						 "101001010001010110111110",
						 "101001010001011000100110",
						 "101001010001011010001110",
						 "101001010001011011110110",
						 "101001010001011101011110",
						 "101001010001011111000110",
						 "101001010001100000101110",
						 "101001010001100010010110",
						 "101001010001100011111110",
						 "101001010001100101100110",
						 "101001010001100111001110",
						 "101001010001101000110110",
						 "101001010001101010011110",
						 "101001010001101100000110",
						 "101001010001010011101110",
						 "101001010001010101010101",
						 "101001010001010110111100",
						 "101001010001011000100011",
						 "101001010001011010001010",
						 "101001010001011011110001",
						 "101001010001011101011000",
						 "101001010001011110111111",
						 "101001010001100000100110",
						 "101001010001100010001101",
						 "101001010001100011110100",
						 "101001010001100101011011",
						 "101001010001100111000010",
						 "101001010001101000101001",
						 "101001010001101010010000",
						 "101001010001101011110111",
						 "101001010001010011101110",
						 "101001010001010101010101",
						 "101001010001010110111100",
						 "101001010001011000100011",
						 "101001010001011010001010",
						 "101001010001011011110001",
						 "101001010001011101011000",
						 "101001010001011110111111",
						 "101001010001100000100110",
						 "101001010001100010001101",
						 "101001010001100011110100",
						 "101001010001100101011011",
						 "101001010001100111000010",
						 "101001010001101000101001",
						 "101001010001101010010000",
						 "101001010001101011110111",
						 "101001010001010011101110",
						 "101001010001010101010100",
						 "101001010001010110111010",
						 "101001010001011000100000",
						 "101001010001011010000110",
						 "101001010001011011101100",
						 "101001010001011101010010",
						 "101001010001011110111000",
						 "101001010001100000011110",
						 "101001010001100010000100",
						 "101001010001100011101010",
						 "101001010001100101010000",
						 "101001010001100110110110",
						 "101001010001101000011100",
						 "101001010001101010000010",
						 "101001010001101011101000",
						 "101001010011110110101100",
						 "101001010011111000010010",
						 "101001010011111001111000",
						 "101001010011111011011110",
						 "101001010011111101000100",
						 "101001010011111110101010",
						 "101001010100000000010000",
						 "101001010100000001110110",
						 "101001010100000011011100",
						 "101001010100000101000010",
						 "101001010100000110101000",
						 "101001010100001000001110",
						 "101001010100001001110100",
						 "101001010100001011011010",
						 "101001010100001101000000",
						 "101001010100001110100110",
						 "101001010011110110101100",
						 "101001010011111000010010",
						 "101001010011111001111000",
						 "101001010011111011011110",
						 "101001010011111101000100",
						 "101001010011111110101010",
						 "101001010100000000010000",
						 "101001010100000001110110",
						 "101001010100000011011100",
						 "101001010100000101000010",
						 "101001010100000110101000",
						 "101001010100001000001110",
						 "101001010100001001110100",
						 "101001010100001011011010",
						 "101001010100001101000000",
						 "101001010100001110100110",
						 "101001010011110110101100",
						 "101001010011111000010001",
						 "101001010011111001110110",
						 "101001010011111011011011",
						 "101001010011111101000000",
						 "101001010011111110100101",
						 "101001010100000000001010",
						 "101001010100000001101111",
						 "101001010100000011010100",
						 "101001010100000100111001",
						 "101001010100000110011110",
						 "101001010100001000000011",
						 "101001010100001001101000",
						 "101001010100001011001101",
						 "101001010100001100110010",
						 "101001010100001110010111",
						 "101001010011110110101100",
						 "101001010011111000010001",
						 "101001010011111001110110",
						 "101001010011111011011011",
						 "101001010011111101000000",
						 "101001010011111110100101",
						 "101001010100000000001010",
						 "101001010100000001101111",
						 "101001010100000011010100",
						 "101001010100000100111001",
						 "101001010100000110011110",
						 "101001010100001000000011",
						 "101001010100001001101000",
						 "101001010100001011001101",
						 "101001010100001100110010",
						 "101001010100001110010111",
						 "101001010011110110101100",
						 "101001010011111000010001",
						 "101001010011111001110110",
						 "101001010011111011011011",
						 "101001010011111101000000",
						 "101001010011111110100101",
						 "101001010100000000001010",
						 "101001010100000001101111",
						 "101001010100000011010100",
						 "101001010100000100111001",
						 "101001010100000110011110",
						 "101001010100001000000011",
						 "101001010100001001101000",
						 "101001010100001011001101",
						 "101001010100001100110010",
						 "101001010100001110010111",
						 "101001010011110110101100",
						 "101001010011111000010000",
						 "101001010011111001110100",
						 "101001010011111011011000",
						 "101001010011111100111100",
						 "101001010011111110100000",
						 "101001010100000000000100",
						 "101001010100000001101000",
						 "101001010100000011001100",
						 "101001010100000100110000",
						 "101001010100000110010100",
						 "101001010100000111111000",
						 "101001010100001001011100",
						 "101001010100001011000000",
						 "101001010100001100100100",
						 "101001010100001110001000",
						 "101001010110011001101010",
						 "101001010110011011001110",
						 "101001010110011100110010",
						 "101001010110011110010110",
						 "101001010110011111111010",
						 "101001010110100001011110",
						 "101001010110100011000010",
						 "101001010110100100100110",
						 "101001010110100110001010",
						 "101001010110100111101110",
						 "101001010110101001010010",
						 "101001010110101010110110",
						 "101001010110101100011010",
						 "101001010110101101111110",
						 "101001010110101111100010",
						 "101001010110110001000110",
						 "101001010110011001101010",
						 "101001010110011011001110",
						 "101001010110011100110010",
						 "101001010110011110010110",
						 "101001010110011111111010",
						 "101001010110100001011110",
						 "101001010110100011000010",
						 "101001010110100100100110",
						 "101001010110100110001010",
						 "101001010110100111101110",
						 "101001010110101001010010",
						 "101001010110101010110110",
						 "101001010110101100011010",
						 "101001010110101101111110",
						 "101001010110101111100010",
						 "101001010110110001000110",
						 "101001010110011001101010",
						 "101001010110011011001101",
						 "101001010110011100110000",
						 "101001010110011110010011",
						 "101001010110011111110110",
						 "101001010110100001011001",
						 "101001010110100010111100",
						 "101001010110100100011111",
						 "101001010110100110000010",
						 "101001010110100111100101",
						 "101001010110101001001000",
						 "101001010110101010101011",
						 "101001010110101100001110",
						 "101001010110101101110001",
						 "101001010110101111010100",
						 "101001010110110000110111",
						 "101001010110011001101010",
						 "101001010110011011001101",
						 "101001010110011100110000",
						 "101001010110011110010011",
						 "101001010110011111110110",
						 "101001010110100001011001",
						 "101001010110100010111100",
						 "101001010110100100011111",
						 "101001010110100110000010",
						 "101001010110100111100101",
						 "101001010110101001001000",
						 "101001010110101010101011",
						 "101001010110101100001110",
						 "101001010110101101110001",
						 "101001010110101111010100",
						 "101001010110110000110111",
						 "101001010110011001101010",
						 "101001010110011011001100",
						 "101001010110011100101110",
						 "101001010110011110010000",
						 "101001010110011111110010",
						 "101001010110100001010100",
						 "101001010110100010110110",
						 "101001010110100100011000",
						 "101001010110100101111010",
						 "101001010110100111011100",
						 "101001010110101000111110",
						 "101001010110101010100000",
						 "101001010110101100000010",
						 "101001010110101101100100",
						 "101001010110101111000110",
						 "101001010110110000101000",
						 "101001010110011001101010",
						 "101001010110011011001100",
						 "101001010110011100101110",
						 "101001010110011110010000",
						 "101001010110011111110010",
						 "101001010110100001010100",
						 "101001010110100010110110",
						 "101001010110100100011000",
						 "101001010110100101111010",
						 "101001010110100111011100",
						 "101001010110101000111110",
						 "101001010110101010100000",
						 "101001010110101100000010",
						 "101001010110101101100100",
						 "101001010110101111000110",
						 "101001010110110000101000",
						 "101001010110011001101010",
						 "101001010110011011001100",
						 "101001010110011100101110",
						 "101001010110011110010000",
						 "101001010110011111110010",
						 "101001010110100001010100",
						 "101001010110100010110110",
						 "101001010110100100011000",
						 "101001010110100101111010",
						 "101001010110100111011100",
						 "101001010110101000111110",
						 "101001010110101010100000",
						 "101001010110101100000010",
						 "101001010110101101100100",
						 "101001010110101111000110",
						 "101001010110110000101000",
						 "101001011000111100101000",
						 "101001011000111110001001",
						 "101001011000111111101010",
						 "101001011001000001001011",
						 "101001011001000010101100",
						 "101001011001000100001101",
						 "101001011001000101101110",
						 "101001011001000111001111",
						 "101001011001001000110000",
						 "101001011001001010010001",
						 "101001011001001011110010",
						 "101001011001001101010011",
						 "101001011001001110110100",
						 "101001011001010000010101",
						 "101001011001010001110110",
						 "101001011001010011010111",
						 "101001011000111100101000",
						 "101001011000111110001001",
						 "101001011000111111101010",
						 "101001011001000001001011",
						 "101001011001000010101100",
						 "101001011001000100001101",
						 "101001011001000101101110",
						 "101001011001000111001111",
						 "101001011001001000110000",
						 "101001011001001010010001",
						 "101001011001001011110010",
						 "101001011001001101010011",
						 "101001011001001110110100",
						 "101001011001010000010101",
						 "101001011001010001110110",
						 "101001011001010011010111",
						 "101001011000111100101000",
						 "101001011000111110001001",
						 "101001011000111111101010",
						 "101001011001000001001011",
						 "101001011001000010101100",
						 "101001011001000100001101",
						 "101001011001000101101110",
						 "101001011001000111001111",
						 "101001011001001000110000",
						 "101001011001001010010001",
						 "101001011001001011110010",
						 "101001011001001101010011",
						 "101001011001001110110100",
						 "101001011001010000010101",
						 "101001011001010001110110",
						 "101001011001010011010111",
						 "101001011000111100101000",
						 "101001011000111110001000",
						 "101001011000111111101000",
						 "101001011001000001001000",
						 "101001011001000010101000",
						 "101001011001000100001000",
						 "101001011001000101101000",
						 "101001011001000111001000",
						 "101001011001001000101000",
						 "101001011001001010001000",
						 "101001011001001011101000",
						 "101001011001001101001000",
						 "101001011001001110101000",
						 "101001011001010000001000",
						 "101001011001010001101000",
						 "101001011001010011001000",
						 "101001011000111100101000",
						 "101001011000111110001000",
						 "101001011000111111101000",
						 "101001011001000001001000",
						 "101001011001000010101000",
						 "101001011001000100001000",
						 "101001011001000101101000",
						 "101001011001000111001000",
						 "101001011001001000101000",
						 "101001011001001010001000",
						 "101001011001001011101000",
						 "101001011001001101001000",
						 "101001011001001110101000",
						 "101001011001010000001000",
						 "101001011001010001101000",
						 "101001011001010011001000",
						 "101001011000111100101000",
						 "101001011000111110001000",
						 "101001011000111111101000",
						 "101001011001000001001000",
						 "101001011001000010101000",
						 "101001011001000100001000",
						 "101001011001000101101000",
						 "101001011001000111001000",
						 "101001011001001000101000",
						 "101001011001001010001000",
						 "101001011001001011101000",
						 "101001011001001101001000",
						 "101001011001001110101000",
						 "101001011001010000001000",
						 "101001011001010001101000",
						 "101001011001010011001000",
						 "101001011000111100101000",
						 "101001011000111110000111",
						 "101001011000111111100110",
						 "101001011001000001000101",
						 "101001011001000010100100",
						 "101001011001000100000011",
						 "101001011001000101100010",
						 "101001011001000111000001",
						 "101001011001001000100000",
						 "101001011001001001111111",
						 "101001011001001011011110",
						 "101001011001001100111101",
						 "101001011001001110011100",
						 "101001011001001111111011",
						 "101001011001010001011010",
						 "101001011001010010111001",
						 "101001011011011111100110",
						 "101001011011100001000101",
						 "101001011011100010100100",
						 "101001011011100100000011",
						 "101001011011100101100010",
						 "101001011011100111000001",
						 "101001011011101000100000",
						 "101001011011101001111111",
						 "101001011011101011011110",
						 "101001011011101100111101",
						 "101001011011101110011100",
						 "101001011011101111111011",
						 "101001011011110001011010",
						 "101001011011110010111001",
						 "101001011011110100011000",
						 "101001011011110101110111",
						 "101001011011011111100110",
						 "101001011011100001000100",
						 "101001011011100010100010",
						 "101001011011100100000000",
						 "101001011011100101011110",
						 "101001011011100110111100",
						 "101001011011101000011010",
						 "101001011011101001111000",
						 "101001011011101011010110",
						 "101001011011101100110100",
						 "101001011011101110010010",
						 "101001011011101111110000",
						 "101001011011110001001110",
						 "101001011011110010101100",
						 "101001011011110100001010",
						 "101001011011110101101000",
						 "101001011011011111100110",
						 "101001011011100001000100",
						 "101001011011100010100010",
						 "101001011011100100000000",
						 "101001011011100101011110",
						 "101001011011100110111100",
						 "101001011011101000011010",
						 "101001011011101001111000",
						 "101001011011101011010110",
						 "101001011011101100110100",
						 "101001011011101110010010",
						 "101001011011101111110000",
						 "101001011011110001001110",
						 "101001011011110010101100",
						 "101001011011110100001010",
						 "101001011011110101101000",
						 "101001011011011111100110",
						 "101001011011100001000100",
						 "101001011011100010100010",
						 "101001011011100100000000",
						 "101001011011100101011110",
						 "101001011011100110111100",
						 "101001011011101000011010",
						 "101001011011101001111000",
						 "101001011011101011010110",
						 "101001011011101100110100",
						 "101001011011101110010010",
						 "101001011011101111110000",
						 "101001011011110001001110",
						 "101001011011110010101100",
						 "101001011011110100001010",
						 "101001011011110101101000",
						 "101001011011011111100110",
						 "101001011011100001000011",
						 "101001011011100010100000",
						 "101001011011100011111101",
						 "101001011011100101011010",
						 "101001011011100110110111",
						 "101001011011101000010100",
						 "101001011011101001110001",
						 "101001011011101011001110",
						 "101001011011101100101011",
						 "101001011011101110001000",
						 "101001011011101111100101",
						 "101001011011110001000010",
						 "101001011011110010011111",
						 "101001011011110011111100",
						 "101001011011110101011001",
						 "101001011011011111100110",
						 "101001011011100001000011",
						 "101001011011100010100000",
						 "101001011011100011111101",
						 "101001011011100101011010",
						 "101001011011100110110111",
						 "101001011011101000010100",
						 "101001011011101001110001",
						 "101001011011101011001110",
						 "101001011011101100101011",
						 "101001011011101110001000",
						 "101001011011101111100101",
						 "101001011011110001000010",
						 "101001011011110010011111",
						 "101001011011110011111100",
						 "101001011011110101011001",
						 "101001011011011111100110",
						 "101001011011100001000011",
						 "101001011011100010100000",
						 "101001011011100011111101",
						 "101001011011100101011010",
						 "101001011011100110110111",
						 "101001011011101000010100",
						 "101001011011101001110001",
						 "101001011011101011001110",
						 "101001011011101100101011",
						 "101001011011101110001000",
						 "101001011011101111100101",
						 "101001011011110001000010",
						 "101001011011110010011111",
						 "101001011011110011111100",
						 "101001011011110101011001",
						 "101001011110000010100100",
						 "101001011110000100000000",
						 "101001011110000101011100",
						 "101001011110000110111000",
						 "101001011110001000010100",
						 "101001011110001001110000",
						 "101001011110001011001100",
						 "101001011110001100101000",
						 "101001011110001110000100",
						 "101001011110001111100000",
						 "101001011110010000111100",
						 "101001011110010010011000",
						 "101001011110010011110100",
						 "101001011110010101010000",
						 "101001011110010110101100",
						 "101001011110011000001000",
						 "101001011110000010100100",
						 "101001011110000100000000",
						 "101001011110000101011100",
						 "101001011110000110111000",
						 "101001011110001000010100",
						 "101001011110001001110000",
						 "101001011110001011001100",
						 "101001011110001100101000",
						 "101001011110001110000100",
						 "101001011110001111100000",
						 "101001011110010000111100",
						 "101001011110010010011000",
						 "101001011110010011110100",
						 "101001011110010101010000",
						 "101001011110010110101100",
						 "101001011110011000001000",
						 "101001011110000010100100",
						 "101001011110000100000000",
						 "101001011110000101011100",
						 "101001011110000110111000",
						 "101001011110001000010100",
						 "101001011110001001110000",
						 "101001011110001011001100",
						 "101001011110001100101000",
						 "101001011110001110000100",
						 "101001011110001111100000",
						 "101001011110010000111100",
						 "101001011110010010011000",
						 "101001011110010011110100",
						 "101001011110010101010000",
						 "101001011110010110101100",
						 "101001011110011000001000",
						 "101001011110000010100100",
						 "101001011110000011111111",
						 "101001011110000101011010",
						 "101001011110000110110101",
						 "101001011110001000010000",
						 "101001011110001001101011",
						 "101001011110001011000110",
						 "101001011110001100100001",
						 "101001011110001101111100",
						 "101001011110001111010111",
						 "101001011110010000110010",
						 "101001011110010010001101",
						 "101001011110010011101000",
						 "101001011110010101000011",
						 "101001011110010110011110",
						 "101001011110010111111001",
						 "101001011110000010100100",
						 "101001011110000011111111",
						 "101001011110000101011010",
						 "101001011110000110110101",
						 "101001011110001000010000",
						 "101001011110001001101011",
						 "101001011110001011000110",
						 "101001011110001100100001",
						 "101001011110001101111100",
						 "101001011110001111010111",
						 "101001011110010000110010",
						 "101001011110010010001101",
						 "101001011110010011101000",
						 "101001011110010101000011",
						 "101001011110010110011110",
						 "101001011110010111111001",
						 "101001011110000010100100",
						 "101001011110000011111110",
						 "101001011110000101011000",
						 "101001011110000110110010",
						 "101001011110001000001100",
						 "101001011110001001100110",
						 "101001011110001011000000",
						 "101001011110001100011010",
						 "101001011110001101110100",
						 "101001011110001111001110",
						 "101001011110010000101000",
						 "101001011110010010000010",
						 "101001011110010011011100",
						 "101001011110010100110110",
						 "101001011110010110010000",
						 "101001011110010111101010",
						 "101001011110000010100100",
						 "101001011110000011111110",
						 "101001011110000101011000",
						 "101001011110000110110010",
						 "101001011110001000001100",
						 "101001011110001001100110",
						 "101001011110001011000000",
						 "101001011110001100011010",
						 "101001011110001101110100",
						 "101001011110001111001110",
						 "101001011110010000101000",
						 "101001011110010010000010",
						 "101001011110010011011100",
						 "101001011110010100110110",
						 "101001011110010110010000",
						 "101001011110010111101010",
						 "101001100000100101100010",
						 "101001100000100110111100",
						 "101001100000101000010110",
						 "101001100000101001110000",
						 "101001100000101011001010",
						 "101001100000101100100100",
						 "101001100000101101111110",
						 "101001100000101111011000",
						 "101001100000110000110010",
						 "101001100000110010001100",
						 "101001100000110011100110",
						 "101001100000110101000000",
						 "101001100000110110011010",
						 "101001100000110111110100",
						 "101001100000111001001110",
						 "101001100000111010101000",
						 "101001100000100101100010",
						 "101001100000100110111011",
						 "101001100000101000010100",
						 "101001100000101001101101",
						 "101001100000101011000110",
						 "101001100000101100011111",
						 "101001100000101101111000",
						 "101001100000101111010001",
						 "101001100000110000101010",
						 "101001100000110010000011",
						 "101001100000110011011100",
						 "101001100000110100110101",
						 "101001100000110110001110",
						 "101001100000110111100111",
						 "101001100000111001000000",
						 "101001100000111010011001",
						 "101001100000100101100010",
						 "101001100000100110111011",
						 "101001100000101000010100",
						 "101001100000101001101101",
						 "101001100000101011000110",
						 "101001100000101100011111",
						 "101001100000101101111000",
						 "101001100000101111010001",
						 "101001100000110000101010",
						 "101001100000110010000011",
						 "101001100000110011011100",
						 "101001100000110100110101",
						 "101001100000110110001110",
						 "101001100000110111100111",
						 "101001100000111001000000",
						 "101001100000111010011001",
						 "101001100000100101100010",
						 "101001100000100110111011",
						 "101001100000101000010100",
						 "101001100000101001101101",
						 "101001100000101011000110",
						 "101001100000101100011111",
						 "101001100000101101111000",
						 "101001100000101111010001",
						 "101001100000110000101010",
						 "101001100000110010000011",
						 "101001100000110011011100",
						 "101001100000110100110101",
						 "101001100000110110001110",
						 "101001100000110111100111",
						 "101001100000111001000000",
						 "101001100000111010011001",
						 "101001100000100101100010",
						 "101001100000100110111010",
						 "101001100000101000010010",
						 "101001100000101001101010",
						 "101001100000101011000010",
						 "101001100000101100011010",
						 "101001100000101101110010",
						 "101001100000101111001010",
						 "101001100000110000100010",
						 "101001100000110001111010",
						 "101001100000110011010010",
						 "101001100000110100101010",
						 "101001100000110110000010",
						 "101001100000110111011010",
						 "101001100000111000110010",
						 "101001100000111010001010",
						 "101001100000100101100010",
						 "101001100000100110111010",
						 "101001100000101000010010",
						 "101001100000101001101010",
						 "101001100000101011000010",
						 "101001100000101100011010",
						 "101001100000101101110010",
						 "101001100000101111001010",
						 "101001100000110000100010",
						 "101001100000110001111010",
						 "101001100000110011010010",
						 "101001100000110100101010",
						 "101001100000110110000010",
						 "101001100000110111011010",
						 "101001100000111000110010",
						 "101001100000111010001010",
						 "101001100000100101100010",
						 "101001100000100110111010",
						 "101001100000101000010010",
						 "101001100000101001101010",
						 "101001100000101011000010",
						 "101001100000101100011010",
						 "101001100000101101110010",
						 "101001100000101111001010",
						 "101001100000110000100010",
						 "101001100000110001111010",
						 "101001100000110011010010",
						 "101001100000110100101010",
						 "101001100000110110000010",
						 "101001100000110111011010",
						 "101001100000111000110010",
						 "101001100000111010001010",
						 "101001100011001000100000",
						 "101001100011001001110111",
						 "101001100011001011001110",
						 "101001100011001100100101",
						 "101001100011001101111100",
						 "101001100011001111010011",
						 "101001100011010000101010",
						 "101001100011010010000001",
						 "101001100011010011011000",
						 "101001100011010100101111",
						 "101001100011010110000110",
						 "101001100011010111011101",
						 "101001100011011000110100",
						 "101001100011011010001011",
						 "101001100011011011100010",
						 "101001100011011100111001",
						 "101001100011001000100000",
						 "101001100011001001110111",
						 "101001100011001011001110",
						 "101001100011001100100101",
						 "101001100011001101111100",
						 "101001100011001111010011",
						 "101001100011010000101010",
						 "101001100011010010000001",
						 "101001100011010011011000",
						 "101001100011010100101111",
						 "101001100011010110000110",
						 "101001100011010111011101",
						 "101001100011011000110100",
						 "101001100011011010001011",
						 "101001100011011011100010",
						 "101001100011011100111001",
						 "101001100011001000100000",
						 "101001100011001001110110",
						 "101001100011001011001100",
						 "101001100011001100100010",
						 "101001100011001101111000",
						 "101001100011001111001110",
						 "101001100011010000100100",
						 "101001100011010001111010",
						 "101001100011010011010000",
						 "101001100011010100100110",
						 "101001100011010101111100",
						 "101001100011010111010010",
						 "101001100011011000101000",
						 "101001100011011001111110",
						 "101001100011011011010100",
						 "101001100011011100101010",
						 "101001100011001000100000",
						 "101001100011001001110110",
						 "101001100011001011001100",
						 "101001100011001100100010",
						 "101001100011001101111000",
						 "101001100011001111001110",
						 "101001100011010000100100",
						 "101001100011010001111010",
						 "101001100011010011010000",
						 "101001100011010100100110",
						 "101001100011010101111100",
						 "101001100011010111010010",
						 "101001100011011000101000",
						 "101001100011011001111110",
						 "101001100011011011010100",
						 "101001100011011100101010",
						 "101001100011001000100000",
						 "101001100011001001110110",
						 "101001100011001011001100",
						 "101001100011001100100010",
						 "101001100011001101111000",
						 "101001100011001111001110",
						 "101001100011010000100100",
						 "101001100011010001111010",
						 "101001100011010011010000",
						 "101001100011010100100110",
						 "101001100011010101111100",
						 "101001100011010111010010",
						 "101001100011011000101000",
						 "101001100011011001111110",
						 "101001100011011011010100",
						 "101001100011011100101010",
						 "101001100011001000100000",
						 "101001100011001001110101",
						 "101001100011001011001010",
						 "101001100011001100011111",
						 "101001100011001101110100",
						 "101001100011001111001001",
						 "101001100011010000011110",
						 "101001100011010001110011",
						 "101001100011010011001000",
						 "101001100011010100011101",
						 "101001100011010101110010",
						 "101001100011010111000111",
						 "101001100011011000011100",
						 "101001100011011001110001",
						 "101001100011011011000110",
						 "101001100011011100011011",
						 "101001100011001000100000",
						 "101001100011001001110101",
						 "101001100011001011001010",
						 "101001100011001100011111",
						 "101001100011001101110100",
						 "101001100011001111001001",
						 "101001100011010000011110",
						 "101001100011010001110011",
						 "101001100011010011001000",
						 "101001100011010100011101",
						 "101001100011010101110010",
						 "101001100011010111000111",
						 "101001100011011000011100",
						 "101001100011011001110001",
						 "101001100011011011000110",
						 "101001100011011100011011",
						 "101001100011001000100000",
						 "101001100011001001110101",
						 "101001100011001011001010",
						 "101001100011001100011111",
						 "101001100011001101110100",
						 "101001100011001111001001",
						 "101001100011010000011110",
						 "101001100011010001110011",
						 "101001100011010011001000",
						 "101001100011010100011101",
						 "101001100011010101110010",
						 "101001100011010111000111",
						 "101001100011011000011100",
						 "101001100011011001110001",
						 "101001100011011011000110",
						 "101001100011011100011011",
						 "101001100101101011011110",
						 "101001100101101100110010",
						 "101001100101101110000110",
						 "101001100101101111011010",
						 "101001100101110000101110",
						 "101001100101110010000010",
						 "101001100101110011010110",
						 "101001100101110100101010",
						 "101001100101110101111110",
						 "101001100101110111010010",
						 "101001100101111000100110",
						 "101001100101111001111010",
						 "101001100101111011001110",
						 "101001100101111100100010",
						 "101001100101111101110110",
						 "101001100101111111001010",
						 "101001100101101011011110",
						 "101001100101101100110010",
						 "101001100101101110000110",
						 "101001100101101111011010",
						 "101001100101110000101110",
						 "101001100101110010000010",
						 "101001100101110011010110",
						 "101001100101110100101010",
						 "101001100101110101111110",
						 "101001100101110111010010",
						 "101001100101111000100110",
						 "101001100101111001111010",
						 "101001100101111011001110",
						 "101001100101111100100010",
						 "101001100101111101110110",
						 "101001100101111111001010",
						 "101001100101101011011110",
						 "101001100101101100110001",
						 "101001100101101110000100",
						 "101001100101101111010111",
						 "101001100101110000101010",
						 "101001100101110001111101",
						 "101001100101110011010000",
						 "101001100101110100100011",
						 "101001100101110101110110",
						 "101001100101110111001001",
						 "101001100101111000011100",
						 "101001100101111001101111",
						 "101001100101111011000010",
						 "101001100101111100010101",
						 "101001100101111101101000",
						 "101001100101111110111011",
						 "101001100101101011011110",
						 "101001100101101100110001",
						 "101001100101101110000100",
						 "101001100101101111010111",
						 "101001100101110000101010",
						 "101001100101110001111101",
						 "101001100101110011010000",
						 "101001100101110100100011",
						 "101001100101110101110110",
						 "101001100101110111001001",
						 "101001100101111000011100",
						 "101001100101111001101111",
						 "101001100101111011000010",
						 "101001100101111100010101",
						 "101001100101111101101000",
						 "101001100101111110111011",
						 "101001100101101011011110",
						 "101001100101101100110001",
						 "101001100101101110000100",
						 "101001100101101111010111",
						 "101001100101110000101010",
						 "101001100101110001111101",
						 "101001100101110011010000",
						 "101001100101110100100011",
						 "101001100101110101110110",
						 "101001100101110111001001",
						 "101001100101111000011100",
						 "101001100101111001101111",
						 "101001100101111011000010",
						 "101001100101111100010101",
						 "101001100101111101101000",
						 "101001100101111110111011",
						 "101001100101101011011110",
						 "101001100101101100110000",
						 "101001100101101110000010",
						 "101001100101101111010100",
						 "101001100101110000100110",
						 "101001100101110001111000",
						 "101001100101110011001010",
						 "101001100101110100011100",
						 "101001100101110101101110",
						 "101001100101110111000000",
						 "101001100101111000010010",
						 "101001100101111001100100",
						 "101001100101111010110110",
						 "101001100101111100001000",
						 "101001100101111101011010",
						 "101001100101111110101100",
						 "101001100101101011011110",
						 "101001100101101100110000",
						 "101001100101101110000010",
						 "101001100101101111010100",
						 "101001100101110000100110",
						 "101001100101110001111000",
						 "101001100101110011001010",
						 "101001100101110100011100",
						 "101001100101110101101110",
						 "101001100101110111000000",
						 "101001100101111000010010",
						 "101001100101111001100100",
						 "101001100101111010110110",
						 "101001100101111100001000",
						 "101001100101111101011010",
						 "101001100101111110101100",
						 "101001101000001110011100",
						 "101001101000001111101110",
						 "101001101000010001000000",
						 "101001101000010010010010",
						 "101001101000010011100100",
						 "101001101000010100110110",
						 "101001101000010110001000",
						 "101001101000010111011010",
						 "101001101000011000101100",
						 "101001101000011001111110",
						 "101001101000011011010000",
						 "101001101000011100100010",
						 "101001101000011101110100",
						 "101001101000011111000110",
						 "101001101000100000011000",
						 "101001101000100001101010",
						 "101001101000001110011100",
						 "101001101000001111101101",
						 "101001101000010000111110",
						 "101001101000010010001111",
						 "101001101000010011100000",
						 "101001101000010100110001",
						 "101001101000010110000010",
						 "101001101000010111010011",
						 "101001101000011000100100",
						 "101001101000011001110101",
						 "101001101000011011000110",
						 "101001101000011100010111",
						 "101001101000011101101000",
						 "101001101000011110111001",
						 "101001101000100000001010",
						 "101001101000100001011011",
						 "101001101000001110011100",
						 "101001101000001111101101",
						 "101001101000010000111110",
						 "101001101000010010001111",
						 "101001101000010011100000",
						 "101001101000010100110001",
						 "101001101000010110000010",
						 "101001101000010111010011",
						 "101001101000011000100100",
						 "101001101000011001110101",
						 "101001101000011011000110",
						 "101001101000011100010111",
						 "101001101000011101101000",
						 "101001101000011110111001",
						 "101001101000100000001010",
						 "101001101000100001011011",
						 "101001101000001110011100",
						 "101001101000001111101101",
						 "101001101000010000111110",
						 "101001101000010010001111",
						 "101001101000010011100000",
						 "101001101000010100110001",
						 "101001101000010110000010",
						 "101001101000010111010011",
						 "101001101000011000100100",
						 "101001101000011001110101",
						 "101001101000011011000110",
						 "101001101000011100010111",
						 "101001101000011101101000",
						 "101001101000011110111001",
						 "101001101000100000001010",
						 "101001101000100001011011",
						 "101001101000001110011100",
						 "101001101000001111101100",
						 "101001101000010000111100",
						 "101001101000010010001100",
						 "101001101000010011011100",
						 "101001101000010100101100",
						 "101001101000010101111100",
						 "101001101000010111001100",
						 "101001101000011000011100",
						 "101001101000011001101100",
						 "101001101000011010111100",
						 "101001101000011100001100",
						 "101001101000011101011100",
						 "101001101000011110101100",
						 "101001101000011111111100",
						 "101001101000100001001100",
						 "101001101000001110011100",
						 "101001101000001111101100",
						 "101001101000010000111100",
						 "101001101000010010001100",
						 "101001101000010011011100",
						 "101001101000010100101100",
						 "101001101000010101111100",
						 "101001101000010111001100",
						 "101001101000011000011100",
						 "101001101000011001101100",
						 "101001101000011010111100",
						 "101001101000011100001100",
						 "101001101000011101011100",
						 "101001101000011110101100",
						 "101001101000011111111100",
						 "101001101000100001001100",
						 "101001101000001110011100",
						 "101001101000001111101011",
						 "101001101000010000111010",
						 "101001101000010010001001",
						 "101001101000010011011000",
						 "101001101000010100100111",
						 "101001101000010101110110",
						 "101001101000010111000101",
						 "101001101000011000010100",
						 "101001101000011001100011",
						 "101001101000011010110010",
						 "101001101000011100000001",
						 "101001101000011101010000",
						 "101001101000011110011111",
						 "101001101000011111101110",
						 "101001101000100000111101",
						 "101001101000001110011100",
						 "101001101000001111101011",
						 "101001101000010000111010",
						 "101001101000010010001001",
						 "101001101000010011011000",
						 "101001101000010100100111",
						 "101001101000010101110110",
						 "101001101000010111000101",
						 "101001101000011000010100",
						 "101001101000011001100011",
						 "101001101000011010110010",
						 "101001101000011100000001",
						 "101001101000011101010000",
						 "101001101000011110011111",
						 "101001101000011111101110",
						 "101001101000100000111101",
						 "101001101000001110011100",
						 "101001101000001111101011",
						 "101001101000010000111010",
						 "101001101000010010001001",
						 "101001101000010011011000",
						 "101001101000010100100111",
						 "101001101000010101110110",
						 "101001101000010111000101",
						 "101001101000011000010100",
						 "101001101000011001100011",
						 "101001101000011010110010",
						 "101001101000011100000001",
						 "101001101000011101010000",
						 "101001101000011110011111",
						 "101001101000011111101110",
						 "101001101000100000111101",
						 "101001101010110001011010",
						 "101001101010110010101000",
						 "101001101010110011110110",
						 "101001101010110101000100",
						 "101001101010110110010010",
						 "101001101010110111100000",
						 "101001101010111000101110",
						 "101001101010111001111100",
						 "101001101010111011001010",
						 "101001101010111100011000",
						 "101001101010111101100110",
						 "101001101010111110110100",
						 "101001101011000000000010",
						 "101001101011000001010000",
						 "101001101011000010011110",
						 "101001101011000011101100",
						 "101001101010110001011010",
						 "101001101010110010101000",
						 "101001101010110011110110",
						 "101001101010110101000100",
						 "101001101010110110010010",
						 "101001101010110111100000",
						 "101001101010111000101110",
						 "101001101010111001111100",
						 "101001101010111011001010",
						 "101001101010111100011000",
						 "101001101010111101100110",
						 "101001101010111110110100",
						 "101001101011000000000010",
						 "101001101011000001010000",
						 "101001101011000010011110",
						 "101001101011000011101100",
						 "101001101010110001011010",
						 "101001101010110010101000",
						 "101001101010110011110110",
						 "101001101010110101000100",
						 "101001101010110110010010",
						 "101001101010110111100000",
						 "101001101010111000101110",
						 "101001101010111001111100",
						 "101001101010111011001010",
						 "101001101010111100011000",
						 "101001101010111101100110",
						 "101001101010111110110100",
						 "101001101011000000000010",
						 "101001101011000001010000",
						 "101001101011000010011110",
						 "101001101011000011101100",
						 "101001101010110001011010",
						 "101001101010110010100111",
						 "101001101010110011110100",
						 "101001101010110101000001",
						 "101001101010110110001110",
						 "101001101010110111011011",
						 "101001101010111000101000",
						 "101001101010111001110101",
						 "101001101010111011000010",
						 "101001101010111100001111",
						 "101001101010111101011100",
						 "101001101010111110101001",
						 "101001101010111111110110",
						 "101001101011000001000011",
						 "101001101011000010010000",
						 "101001101011000011011101",
						 "101001101010110001011010",
						 "101001101010110010100111",
						 "101001101010110011110100",
						 "101001101010110101000001",
						 "101001101010110110001110",
						 "101001101010110111011011",
						 "101001101010111000101000",
						 "101001101010111001110101",
						 "101001101010111011000010",
						 "101001101010111100001111",
						 "101001101010111101011100",
						 "101001101010111110101001",
						 "101001101010111111110110",
						 "101001101011000001000011",
						 "101001101011000010010000",
						 "101001101011000011011101",
						 "101001101010110001011010",
						 "101001101010110010100110",
						 "101001101010110011110010",
						 "101001101010110100111110",
						 "101001101010110110001010",
						 "101001101010110111010110",
						 "101001101010111000100010",
						 "101001101010111001101110",
						 "101001101010111010111010",
						 "101001101010111100000110",
						 "101001101010111101010010",
						 "101001101010111110011110",
						 "101001101010111111101010",
						 "101001101011000000110110",
						 "101001101011000010000010",
						 "101001101011000011001110",
						 "101001101010110001011010",
						 "101001101010110010100110",
						 "101001101010110011110010",
						 "101001101010110100111110",
						 "101001101010110110001010",
						 "101001101010110111010110",
						 "101001101010111000100010",
						 "101001101010111001101110",
						 "101001101010111010111010",
						 "101001101010111100000110",
						 "101001101010111101010010",
						 "101001101010111110011110",
						 "101001101010111111101010",
						 "101001101011000000110110",
						 "101001101011000010000010",
						 "101001101011000011001110",
						 "101001101010110001011010",
						 "101001101010110010100110",
						 "101001101010110011110010",
						 "101001101010110100111110",
						 "101001101010110110001010",
						 "101001101010110111010110",
						 "101001101010111000100010",
						 "101001101010111001101110",
						 "101001101010111010111010",
						 "101001101010111100000110",
						 "101001101010111101010010",
						 "101001101010111110011110",
						 "101001101010111111101010",
						 "101001101011000000110110",
						 "101001101011000010000010",
						 "101001101011000011001110",
						 "101001101101010100011000",
						 "101001101101010101100011",
						 "101001101101010110101110",
						 "101001101101010111111001",
						 "101001101101011001000100",
						 "101001101101011010001111",
						 "101001101101011011011010",
						 "101001101101011100100101",
						 "101001101101011101110000",
						 "101001101101011110111011",
						 "101001101101100000000110",
						 "101001101101100001010001",
						 "101001101101100010011100",
						 "101001101101100011100111",
						 "101001101101100100110010",
						 "101001101101100101111101",
						 "101001101101010100011000",
						 "101001101101010101100011",
						 "101001101101010110101110",
						 "101001101101010111111001",
						 "101001101101011001000100",
						 "101001101101011010001111",
						 "101001101101011011011010",
						 "101001101101011100100101",
						 "101001101101011101110000",
						 "101001101101011110111011",
						 "101001101101100000000110",
						 "101001101101100001010001",
						 "101001101101100010011100",
						 "101001101101100011100111",
						 "101001101101100100110010",
						 "101001101101100101111101",
						 "101001101101010100011000",
						 "101001101101010101100011",
						 "101001101101010110101110",
						 "101001101101010111111001",
						 "101001101101011001000100",
						 "101001101101011010001111",
						 "101001101101011011011010",
						 "101001101101011100100101",
						 "101001101101011101110000",
						 "101001101101011110111011",
						 "101001101101100000000110",
						 "101001101101100001010001",
						 "101001101101100010011100",
						 "101001101101100011100111",
						 "101001101101100100110010",
						 "101001101101100101111101",
						 "101001101101010100011000",
						 "101001101101010101100010",
						 "101001101101010110101100",
						 "101001101101010111110110",
						 "101001101101011001000000",
						 "101001101101011010001010",
						 "101001101101011011010100",
						 "101001101101011100011110",
						 "101001101101011101101000",
						 "101001101101011110110010",
						 "101001101101011111111100",
						 "101001101101100001000110",
						 "101001101101100010010000",
						 "101001101101100011011010",
						 "101001101101100100100100",
						 "101001101101100101101110",
						 "101001101101010100011000",
						 "101001101101010101100010",
						 "101001101101010110101100",
						 "101001101101010111110110",
						 "101001101101011001000000",
						 "101001101101011010001010",
						 "101001101101011011010100",
						 "101001101101011100011110",
						 "101001101101011101101000",
						 "101001101101011110110010",
						 "101001101101011111111100",
						 "101001101101100001000110",
						 "101001101101100010010000",
						 "101001101101100011011010",
						 "101001101101100100100100",
						 "101001101101100101101110",
						 "101001101101010100011000",
						 "101001101101010101100001",
						 "101001101101010110101010",
						 "101001101101010111110011",
						 "101001101101011000111100",
						 "101001101101011010000101",
						 "101001101101011011001110",
						 "101001101101011100010111",
						 "101001101101011101100000",
						 "101001101101011110101001",
						 "101001101101011111110010",
						 "101001101101100000111011",
						 "101001101101100010000100",
						 "101001101101100011001101",
						 "101001101101100100010110",
						 "101001101101100101011111",
						 "101001101101010100011000",
						 "101001101101010101100001",
						 "101001101101010110101010",
						 "101001101101010111110011",
						 "101001101101011000111100",
						 "101001101101011010000101",
						 "101001101101011011001110",
						 "101001101101011100010111",
						 "101001101101011101100000",
						 "101001101101011110101001",
						 "101001101101011111110010",
						 "101001101101100000111011",
						 "101001101101100010000100",
						 "101001101101100011001101",
						 "101001101101100100010110",
						 "101001101101100101011111",
						 "101001101101010100011000",
						 "101001101101010101100001",
						 "101001101101010110101010",
						 "101001101101010111110011",
						 "101001101101011000111100",
						 "101001101101011010000101",
						 "101001101101011011001110",
						 "101001101101011100010111",
						 "101001101101011101100000",
						 "101001101101011110101001",
						 "101001101101011111110010",
						 "101001101101100000111011",
						 "101001101101100010000100",
						 "101001101101100011001101",
						 "101001101101100100010110",
						 "101001101101100101011111",
						 "101001101101010100011000",
						 "101001101101010101100000",
						 "101001101101010110101000",
						 "101001101101010111110000",
						 "101001101101011000111000",
						 "101001101101011010000000",
						 "101001101101011011001000",
						 "101001101101011100010000",
						 "101001101101011101011000",
						 "101001101101011110100000",
						 "101001101101011111101000",
						 "101001101101100000110000",
						 "101001101101100001111000",
						 "101001101101100011000000",
						 "101001101101100100001000",
						 "101001101101100101010000",
						 "101001101111110111010110",
						 "101001101111111000011110",
						 "101001101111111001100110",
						 "101001101111111010101110",
						 "101001101111111011110110",
						 "101001101111111100111110",
						 "101001101111111110000110",
						 "101001101111111111001110",
						 "101001110000000000010110",
						 "101001110000000001011110",
						 "101001110000000010100110",
						 "101001110000000011101110",
						 "101001110000000100110110",
						 "101001110000000101111110",
						 "101001110000000111000110",
						 "101001110000001000001110",
						 "101001101111110111010110",
						 "101001101111111000011110",
						 "101001101111111001100110",
						 "101001101111111010101110",
						 "101001101111111011110110",
						 "101001101111111100111110",
						 "101001101111111110000110",
						 "101001101111111111001110",
						 "101001110000000000010110",
						 "101001110000000001011110",
						 "101001110000000010100110",
						 "101001110000000011101110",
						 "101001110000000100110110",
						 "101001110000000101111110",
						 "101001110000000111000110",
						 "101001110000001000001110",
						 "101001101111110111010110",
						 "101001101111111000011101",
						 "101001101111111001100100",
						 "101001101111111010101011",
						 "101001101111111011110010",
						 "101001101111111100111001",
						 "101001101111111110000000",
						 "101001101111111111000111",
						 "101001110000000000001110",
						 "101001110000000001010101",
						 "101001110000000010011100",
						 "101001110000000011100011",
						 "101001110000000100101010",
						 "101001110000000101110001",
						 "101001110000000110111000",
						 "101001110000000111111111",
						 "101001101111110111010110",
						 "101001101111111000011101",
						 "101001101111111001100100",
						 "101001101111111010101011",
						 "101001101111111011110010",
						 "101001101111111100111001",
						 "101001101111111110000000",
						 "101001101111111111000111",
						 "101001110000000000001110",
						 "101001110000000001010101",
						 "101001110000000010011100",
						 "101001110000000011100011",
						 "101001110000000100101010",
						 "101001110000000101110001",
						 "101001110000000110111000",
						 "101001110000000111111111",
						 "101001101111110111010110",
						 "101001101111111000011100",
						 "101001101111111001100010",
						 "101001101111111010101000",
						 "101001101111111011101110",
						 "101001101111111100110100",
						 "101001101111111101111010",
						 "101001101111111111000000",
						 "101001110000000000000110",
						 "101001110000000001001100",
						 "101001110000000010010010",
						 "101001110000000011011000",
						 "101001110000000100011110",
						 "101001110000000101100100",
						 "101001110000000110101010",
						 "101001110000000111110000",
						 "101001101111110111010110",
						 "101001101111111000011100",
						 "101001101111111001100010",
						 "101001101111111010101000",
						 "101001101111111011101110",
						 "101001101111111100110100",
						 "101001101111111101111010",
						 "101001101111111111000000",
						 "101001110000000000000110",
						 "101001110000000001001100",
						 "101001110000000010010010",
						 "101001110000000011011000",
						 "101001110000000100011110",
						 "101001110000000101100100",
						 "101001110000000110101010",
						 "101001110000000111110000",
						 "101001101111110111010110",
						 "101001101111111000011100",
						 "101001101111111001100010",
						 "101001101111111010101000",
						 "101001101111111011101110",
						 "101001101111111100110100",
						 "101001101111111101111010",
						 "101001101111111111000000",
						 "101001110000000000000110",
						 "101001110000000001001100",
						 "101001110000000010010010",
						 "101001110000000011011000",
						 "101001110000000100011110",
						 "101001110000000101100100",
						 "101001110000000110101010",
						 "101001110000000111110000",
						 "101001101111110111010110",
						 "101001101111111000011011",
						 "101001101111111001100000",
						 "101001101111111010100101",
						 "101001101111111011101010",
						 "101001101111111100101111",
						 "101001101111111101110100",
						 "101001101111111110111001",
						 "101001101111111111111110",
						 "101001110000000001000011",
						 "101001110000000010001000",
						 "101001110000000011001101",
						 "101001110000000100010010",
						 "101001110000000101010111",
						 "101001110000000110011100",
						 "101001110000000111100001",
						 "101001101111110111010110",
						 "101001101111111000011011",
						 "101001101111111001100000",
						 "101001101111111010100101",
						 "101001101111111011101010",
						 "101001101111111100101111",
						 "101001101111111101110100",
						 "101001101111111110111001",
						 "101001101111111111111110",
						 "101001110000000001000011",
						 "101001110000000010001000",
						 "101001110000000011001101",
						 "101001110000000100010010",
						 "101001110000000101010111",
						 "101001110000000110011100",
						 "101001110000000111100001",
						 "101001110010011010010100",
						 "101001110010011011011001",
						 "101001110010011100011110",
						 "101001110010011101100011",
						 "101001110010011110101000",
						 "101001110010011111101101",
						 "101001110010100000110010",
						 "101001110010100001110111",
						 "101001110010100010111100",
						 "101001110010100100000001",
						 "101001110010100101000110",
						 "101001110010100110001011",
						 "101001110010100111010000",
						 "101001110010101000010101",
						 "101001110010101001011010",
						 "101001110010101010011111",
						 "101001110010011010010100",
						 "101001110010011011011000",
						 "101001110010011100011100",
						 "101001110010011101100000",
						 "101001110010011110100100",
						 "101001110010011111101000",
						 "101001110010100000101100",
						 "101001110010100001110000",
						 "101001110010100010110100",
						 "101001110010100011111000",
						 "101001110010100100111100",
						 "101001110010100110000000",
						 "101001110010100111000100",
						 "101001110010101000001000",
						 "101001110010101001001100",
						 "101001110010101010010000",
						 "101001110010011010010100",
						 "101001110010011011011000",
						 "101001110010011100011100",
						 "101001110010011101100000",
						 "101001110010011110100100",
						 "101001110010011111101000",
						 "101001110010100000101100",
						 "101001110010100001110000",
						 "101001110010100010110100",
						 "101001110010100011111000",
						 "101001110010100100111100",
						 "101001110010100110000000",
						 "101001110010100111000100",
						 "101001110010101000001000",
						 "101001110010101001001100",
						 "101001110010101010010000",
						 "101001110010011010010100",
						 "101001110010011011010111",
						 "101001110010011100011010",
						 "101001110010011101011101",
						 "101001110010011110100000",
						 "101001110010011111100011",
						 "101001110010100000100110",
						 "101001110010100001101001",
						 "101001110010100010101100",
						 "101001110010100011101111",
						 "101001110010100100110010",
						 "101001110010100101110101",
						 "101001110010100110111000",
						 "101001110010100111111011",
						 "101001110010101000111110",
						 "101001110010101010000001",
						 "101001110010011010010100",
						 "101001110010011011010111",
						 "101001110010011100011010",
						 "101001110010011101011101",
						 "101001110010011110100000",
						 "101001110010011111100011",
						 "101001110010100000100110",
						 "101001110010100001101001",
						 "101001110010100010101100",
						 "101001110010100011101111",
						 "101001110010100100110010",
						 "101001110010100101110101",
						 "101001110010100110111000",
						 "101001110010100111111011",
						 "101001110010101000111110",
						 "101001110010101010000001",
						 "101001110010011010010100",
						 "101001110010011011010111",
						 "101001110010011100011010",
						 "101001110010011101011101",
						 "101001110010011110100000",
						 "101001110010011111100011",
						 "101001110010100000100110",
						 "101001110010100001101001",
						 "101001110010100010101100",
						 "101001110010100011101111",
						 "101001110010100100110010",
						 "101001110010100101110101",
						 "101001110010100110111000",
						 "101001110010100111111011",
						 "101001110010101000111110",
						 "101001110010101010000001",
						 "101001110010011010010100",
						 "101001110010011011010110",
						 "101001110010011100011000",
						 "101001110010011101011010",
						 "101001110010011110011100",
						 "101001110010011111011110",
						 "101001110010100000100000",
						 "101001110010100001100010",
						 "101001110010100010100100",
						 "101001110010100011100110",
						 "101001110010100100101000",
						 "101001110010100101101010",
						 "101001110010100110101100",
						 "101001110010100111101110",
						 "101001110010101000110000",
						 "101001110010101001110010",
						 "101001110010011010010100",
						 "101001110010011011010110",
						 "101001110010011100011000",
						 "101001110010011101011010",
						 "101001110010011110011100",
						 "101001110010011111011110",
						 "101001110010100000100000",
						 "101001110010100001100010",
						 "101001110010100010100100",
						 "101001110010100011100110",
						 "101001110010100100101000",
						 "101001110010100101101010",
						 "101001110010100110101100",
						 "101001110010100111101110",
						 "101001110010101000110000",
						 "101001110010101001110010",
						 "101001110010011010010100",
						 "101001110010011011010110",
						 "101001110010011100011000",
						 "101001110010011101011010",
						 "101001110010011110011100",
						 "101001110010011111011110",
						 "101001110010100000100000",
						 "101001110010100001100010",
						 "101001110010100010100100",
						 "101001110010100011100110",
						 "101001110010100100101000",
						 "101001110010100101101010",
						 "101001110010100110101100",
						 "101001110010100111101110",
						 "101001110010101000110000",
						 "101001110010101001110010",
						 "101001110010011010010100",
						 "101001110010011011010101",
						 "101001110010011100010110",
						 "101001110010011101010111",
						 "101001110010011110011000",
						 "101001110010011111011001",
						 "101001110010100000011010",
						 "101001110010100001011011",
						 "101001110010100010011100",
						 "101001110010100011011101",
						 "101001110010100100011110",
						 "101001110010100101011111",
						 "101001110010100110100000",
						 "101001110010100111100001",
						 "101001110010101000100010",
						 "101001110010101001100011",
						 "101001110100111101010010",
						 "101001110100111110010011",
						 "101001110100111111010100",
						 "101001110101000000010101",
						 "101001110101000001010110",
						 "101001110101000010010111",
						 "101001110101000011011000",
						 "101001110101000100011001",
						 "101001110101000101011010",
						 "101001110101000110011011",
						 "101001110101000111011100",
						 "101001110101001000011101",
						 "101001110101001001011110",
						 "101001110101001010011111",
						 "101001110101001011100000",
						 "101001110101001100100001",
						 "101001110100111101010010",
						 "101001110100111110010010",
						 "101001110100111111010010",
						 "101001110101000000010010",
						 "101001110101000001010010",
						 "101001110101000010010010",
						 "101001110101000011010010",
						 "101001110101000100010010",
						 "101001110101000101010010",
						 "101001110101000110010010",
						 "101001110101000111010010",
						 "101001110101001000010010",
						 "101001110101001001010010",
						 "101001110101001010010010",
						 "101001110101001011010010",
						 "101001110101001100010010",
						 "101001110100111101010010",
						 "101001110100111110010010",
						 "101001110100111111010010",
						 "101001110101000000010010",
						 "101001110101000001010010",
						 "101001110101000010010010",
						 "101001110101000011010010",
						 "101001110101000100010010",
						 "101001110101000101010010",
						 "101001110101000110010010",
						 "101001110101000111010010",
						 "101001110101001000010010",
						 "101001110101001001010010",
						 "101001110101001010010010",
						 "101001110101001011010010",
						 "101001110101001100010010",
						 "101001110100111101010010",
						 "101001110100111110010010",
						 "101001110100111111010010",
						 "101001110101000000010010",
						 "101001110101000001010010",
						 "101001110101000010010010",
						 "101001110101000011010010",
						 "101001110101000100010010",
						 "101001110101000101010010",
						 "101001110101000110010010",
						 "101001110101000111010010",
						 "101001110101001000010010",
						 "101001110101001001010010",
						 "101001110101001010010010",
						 "101001110101001011010010",
						 "101001110101001100010010",
						 "101001110100111101010010",
						 "101001110100111110010001",
						 "101001110100111111010000",
						 "101001110101000000001111",
						 "101001110101000001001110",
						 "101001110101000010001101",
						 "101001110101000011001100",
						 "101001110101000100001011",
						 "101001110101000101001010",
						 "101001110101000110001001",
						 "101001110101000111001000",
						 "101001110101001000000111",
						 "101001110101001001000110",
						 "101001110101001010000101",
						 "101001110101001011000100",
						 "101001110101001100000011",
						 "101001110100111101010010",
						 "101001110100111110010001",
						 "101001110100111111010000",
						 "101001110101000000001111",
						 "101001110101000001001110",
						 "101001110101000010001101",
						 "101001110101000011001100",
						 "101001110101000100001011",
						 "101001110101000101001010",
						 "101001110101000110001001",
						 "101001110101000111001000",
						 "101001110101001000000111",
						 "101001110101001001000110",
						 "101001110101001010000101",
						 "101001110101001011000100",
						 "101001110101001100000011",
						 "101001110100111101010010",
						 "101001110100111110010001",
						 "101001110100111111010000",
						 "101001110101000000001111",
						 "101001110101000001001110",
						 "101001110101000010001101",
						 "101001110101000011001100",
						 "101001110101000100001011",
						 "101001110101000101001010",
						 "101001110101000110001001",
						 "101001110101000111001000",
						 "101001110101001000000111",
						 "101001110101001001000110",
						 "101001110101001010000101",
						 "101001110101001011000100",
						 "101001110101001100000011",
						 "101001110100111101010010",
						 "101001110100111110010000",
						 "101001110100111111001110",
						 "101001110101000000001100",
						 "101001110101000001001010",
						 "101001110101000010001000",
						 "101001110101000011000110",
						 "101001110101000100000100",
						 "101001110101000101000010",
						 "101001110101000110000000",
						 "101001110101000110111110",
						 "101001110101000111111100",
						 "101001110101001000111010",
						 "101001110101001001111000",
						 "101001110101001010110110",
						 "101001110101001011110100",
						 "101001110100111101010010",
						 "101001110100111110010000",
						 "101001110100111111001110",
						 "101001110101000000001100",
						 "101001110101000001001010",
						 "101001110101000010001000",
						 "101001110101000011000110",
						 "101001110101000100000100",
						 "101001110101000101000010",
						 "101001110101000110000000",
						 "101001110101000110111110",
						 "101001110101000111111100",
						 "101001110101001000111010",
						 "101001110101001001111000",
						 "101001110101001010110110",
						 "101001110101001011110100",
						 "101001110100111101010010",
						 "101001110100111110001111",
						 "101001110100111111001100",
						 "101001110101000000001001",
						 "101001110101000001000110",
						 "101001110101000010000011",
						 "101001110101000011000000",
						 "101001110101000011111101",
						 "101001110101000100111010",
						 "101001110101000101110111",
						 "101001110101000110110100",
						 "101001110101000111110001",
						 "101001110101001000101110",
						 "101001110101001001101011",
						 "101001110101001010101000",
						 "101001110101001011100101",
						 "101001110111100000010000",
						 "101001110111100001001101",
						 "101001110111100010001010",
						 "101001110111100011000111",
						 "101001110111100100000100",
						 "101001110111100101000001",
						 "101001110111100101111110",
						 "101001110111100110111011",
						 "101001110111100111111000",
						 "101001110111101000110101",
						 "101001110111101001110010",
						 "101001110111101010101111",
						 "101001110111101011101100",
						 "101001110111101100101001",
						 "101001110111101101100110",
						 "101001110111101110100011",
						 "101001110111100000010000",
						 "101001110111100001001101",
						 "101001110111100010001010",
						 "101001110111100011000111",
						 "101001110111100100000100",
						 "101001110111100101000001",
						 "101001110111100101111110",
						 "101001110111100110111011",
						 "101001110111100111111000",
						 "101001110111101000110101",
						 "101001110111101001110010",
						 "101001110111101010101111",
						 "101001110111101011101100",
						 "101001110111101100101001",
						 "101001110111101101100110",
						 "101001110111101110100011",
						 "101001110111100000010000",
						 "101001110111100001001100",
						 "101001110111100010001000",
						 "101001110111100011000100",
						 "101001110111100100000000",
						 "101001110111100100111100",
						 "101001110111100101111000",
						 "101001110111100110110100",
						 "101001110111100111110000",
						 "101001110111101000101100",
						 "101001110111101001101000",
						 "101001110111101010100100",
						 "101001110111101011100000",
						 "101001110111101100011100",
						 "101001110111101101011000",
						 "101001110111101110010100",
						 "101001110111100000010000",
						 "101001110111100001001100",
						 "101001110111100010001000",
						 "101001110111100011000100",
						 "101001110111100100000000",
						 "101001110111100100111100",
						 "101001110111100101111000",
						 "101001110111100110110100",
						 "101001110111100111110000",
						 "101001110111101000101100",
						 "101001110111101001101000",
						 "101001110111101010100100",
						 "101001110111101011100000",
						 "101001110111101100011100",
						 "101001110111101101011000",
						 "101001110111101110010100",
						 "101001110111100000010000",
						 "101001110111100001001011",
						 "101001110111100010000110",
						 "101001110111100011000001",
						 "101001110111100011111100",
						 "101001110111100100110111",
						 "101001110111100101110010",
						 "101001110111100110101101",
						 "101001110111100111101000",
						 "101001110111101000100011",
						 "101001110111101001011110",
						 "101001110111101010011001",
						 "101001110111101011010100",
						 "101001110111101100001111",
						 "101001110111101101001010",
						 "101001110111101110000101",
						 "101001110111100000010000",
						 "101001110111100001001011",
						 "101001110111100010000110",
						 "101001110111100011000001",
						 "101001110111100011111100",
						 "101001110111100100110111",
						 "101001110111100101110010",
						 "101001110111100110101101",
						 "101001110111100111101000",
						 "101001110111101000100011",
						 "101001110111101001011110",
						 "101001110111101010011001",
						 "101001110111101011010100",
						 "101001110111101100001111",
						 "101001110111101101001010",
						 "101001110111101110000101",
						 "101001110111100000010000",
						 "101001110111100001001011",
						 "101001110111100010000110",
						 "101001110111100011000001",
						 "101001110111100011111100",
						 "101001110111100100110111",
						 "101001110111100101110010",
						 "101001110111100110101101",
						 "101001110111100111101000",
						 "101001110111101000100011",
						 "101001110111101001011110",
						 "101001110111101010011001",
						 "101001110111101011010100",
						 "101001110111101100001111",
						 "101001110111101101001010",
						 "101001110111101110000101",
						 "101001110111100000010000",
						 "101001110111100001001010",
						 "101001110111100010000100",
						 "101001110111100010111110",
						 "101001110111100011111000",
						 "101001110111100100110010",
						 "101001110111100101101100",
						 "101001110111100110100110",
						 "101001110111100111100000",
						 "101001110111101000011010",
						 "101001110111101001010100",
						 "101001110111101010001110",
						 "101001110111101011001000",
						 "101001110111101100000010",
						 "101001110111101100111100",
						 "101001110111101101110110",
						 "101001110111100000010000",
						 "101001110111100001001010",
						 "101001110111100010000100",
						 "101001110111100010111110",
						 "101001110111100011111000",
						 "101001110111100100110010",
						 "101001110111100101101100",
						 "101001110111100110100110",
						 "101001110111100111100000",
						 "101001110111101000011010",
						 "101001110111101001010100",
						 "101001110111101010001110",
						 "101001110111101011001000",
						 "101001110111101100000010",
						 "101001110111101100111100",
						 "101001110111101101110110",
						 "101001110111100000010000",
						 "101001110111100001001010",
						 "101001110111100010000100",
						 "101001110111100010111110",
						 "101001110111100011111000",
						 "101001110111100100110010",
						 "101001110111100101101100",
						 "101001110111100110100110",
						 "101001110111100111100000",
						 "101001110111101000011010",
						 "101001110111101001010100",
						 "101001110111101010001110",
						 "101001110111101011001000",
						 "101001110111101100000010",
						 "101001110111101100111100",
						 "101001110111101101110110",
						 "101001110111100000010000",
						 "101001110111100001001001",
						 "101001110111100010000010",
						 "101001110111100010111011",
						 "101001110111100011110100",
						 "101001110111100100101101",
						 "101001110111100101100110",
						 "101001110111100110011111",
						 "101001110111100111011000",
						 "101001110111101000010001",
						 "101001110111101001001010",
						 "101001110111101010000011",
						 "101001110111101010111100",
						 "101001110111101011110101",
						 "101001110111101100101110",
						 "101001110111101101100111",
						 "101001111010000011001110",
						 "101001111010000100000111",
						 "101001111010000101000000",
						 "101001111010000101111001",
						 "101001111010000110110010",
						 "101001111010000111101011",
						 "101001111010001000100100",
						 "101001111010001001011101",
						 "101001111010001010010110",
						 "101001111010001011001111",
						 "101001111010001100001000",
						 "101001111010001101000001",
						 "101001111010001101111010",
						 "101001111010001110110011",
						 "101001111010001111101100",
						 "101001111010010000100101",
						 "101001111010000011001110",
						 "101001111010000100000110",
						 "101001111010000100111110",
						 "101001111010000101110110",
						 "101001111010000110101110",
						 "101001111010000111100110",
						 "101001111010001000011110",
						 "101001111010001001010110",
						 "101001111010001010001110",
						 "101001111010001011000110",
						 "101001111010001011111110",
						 "101001111010001100110110",
						 "101001111010001101101110",
						 "101001111010001110100110",
						 "101001111010001111011110",
						 "101001111010010000010110",
						 "101001111010000011001110",
						 "101001111010000100000110",
						 "101001111010000100111110",
						 "101001111010000101110110",
						 "101001111010000110101110",
						 "101001111010000111100110",
						 "101001111010001000011110",
						 "101001111010001001010110",
						 "101001111010001010001110",
						 "101001111010001011000110",
						 "101001111010001011111110",
						 "101001111010001100110110",
						 "101001111010001101101110",
						 "101001111010001110100110",
						 "101001111010001111011110",
						 "101001111010010000010110",
						 "101001111010000011001110",
						 "101001111010000100000110",
						 "101001111010000100111110",
						 "101001111010000101110110",
						 "101001111010000110101110",
						 "101001111010000111100110",
						 "101001111010001000011110",
						 "101001111010001001010110",
						 "101001111010001010001110",
						 "101001111010001011000110",
						 "101001111010001011111110",
						 "101001111010001100110110",
						 "101001111010001101101110",
						 "101001111010001110100110",
						 "101001111010001111011110",
						 "101001111010010000010110",
						 "101001111010000011001110",
						 "101001111010000100000101",
						 "101001111010000100111100",
						 "101001111010000101110011",
						 "101001111010000110101010",
						 "101001111010000111100001",
						 "101001111010001000011000",
						 "101001111010001001001111",
						 "101001111010001010000110",
						 "101001111010001010111101",
						 "101001111010001011110100",
						 "101001111010001100101011",
						 "101001111010001101100010",
						 "101001111010001110011001",
						 "101001111010001111010000",
						 "101001111010010000000111",
						 "101001111010000011001110",
						 "101001111010000100000101",
						 "101001111010000100111100",
						 "101001111010000101110011",
						 "101001111010000110101010",
						 "101001111010000111100001",
						 "101001111010001000011000",
						 "101001111010001001001111",
						 "101001111010001010000110",
						 "101001111010001010111101",
						 "101001111010001011110100",
						 "101001111010001100101011",
						 "101001111010001101100010",
						 "101001111010001110011001",
						 "101001111010001111010000",
						 "101001111010010000000111",
						 "101001111010000011001110",
						 "101001111010000100000101",
						 "101001111010000100111100",
						 "101001111010000101110011",
						 "101001111010000110101010",
						 "101001111010000111100001",
						 "101001111010001000011000",
						 "101001111010001001001111",
						 "101001111010001010000110",
						 "101001111010001010111101",
						 "101001111010001011110100",
						 "101001111010001100101011",
						 "101001111010001101100010",
						 "101001111010001110011001",
						 "101001111010001111010000",
						 "101001111010010000000111",
						 "101001111010000011001110",
						 "101001111010000100000100",
						 "101001111010000100111010",
						 "101001111010000101110000",
						 "101001111010000110100110",
						 "101001111010000111011100",
						 "101001111010001000010010",
						 "101001111010001001001000",
						 "101001111010001001111110",
						 "101001111010001010110100",
						 "101001111010001011101010",
						 "101001111010001100100000",
						 "101001111010001101010110",
						 "101001111010001110001100",
						 "101001111010001111000010",
						 "101001111010001111111000",
						 "101001111010000011001110",
						 "101001111010000100000100",
						 "101001111010000100111010",
						 "101001111010000101110000",
						 "101001111010000110100110",
						 "101001111010000111011100",
						 "101001111010001000010010",
						 "101001111010001001001000",
						 "101001111010001001111110",
						 "101001111010001010110100",
						 "101001111010001011101010",
						 "101001111010001100100000",
						 "101001111010001101010110",
						 "101001111010001110001100",
						 "101001111010001111000010",
						 "101001111010001111111000",
						 "101001111010000011001110",
						 "101001111010000100000011",
						 "101001111010000100111000",
						 "101001111010000101101101",
						 "101001111010000110100010",
						 "101001111010000111010111",
						 "101001111010001000001100",
						 "101001111010001001000001",
						 "101001111010001001110110",
						 "101001111010001010101011",
						 "101001111010001011100000",
						 "101001111010001100010101",
						 "101001111010001101001010",
						 "101001111010001101111111",
						 "101001111010001110110100",
						 "101001111010001111101001",
						 "101001111010000011001110",
						 "101001111010000100000011",
						 "101001111010000100111000",
						 "101001111010000101101101",
						 "101001111010000110100010",
						 "101001111010000111010111",
						 "101001111010001000001100",
						 "101001111010001001000001",
						 "101001111010001001110110",
						 "101001111010001010101011",
						 "101001111010001011100000",
						 "101001111010001100010101",
						 "101001111010001101001010",
						 "101001111010001101111111",
						 "101001111010001110110100",
						 "101001111010001111101001",
						 "101001111010000011001110",
						 "101001111010000100000011",
						 "101001111010000100111000",
						 "101001111010000101101101",
						 "101001111010000110100010",
						 "101001111010000111010111",
						 "101001111010001000001100",
						 "101001111010001001000001",
						 "101001111010001001110110",
						 "101001111010001010101011",
						 "101001111010001011100000",
						 "101001111010001100010101",
						 "101001111010001101001010",
						 "101001111010001101111111",
						 "101001111010001110110100",
						 "101001111010001111101001",
						 "101001111100100110001100",
						 "101001111100100111000000",
						 "101001111100100111110100",
						 "101001111100101000101000",
						 "101001111100101001011100",
						 "101001111100101010010000",
						 "101001111100101011000100",
						 "101001111100101011111000",
						 "101001111100101100101100",
						 "101001111100101101100000",
						 "101001111100101110010100",
						 "101001111100101111001000",
						 "101001111100101111111100",
						 "101001111100110000110000",
						 "101001111100110001100100",
						 "101001111100110010011000",
						 "101001111100100110001100",
						 "101001111100100111000000",
						 "101001111100100111110100",
						 "101001111100101000101000",
						 "101001111100101001011100",
						 "101001111100101010010000",
						 "101001111100101011000100",
						 "101001111100101011111000",
						 "101001111100101100101100",
						 "101001111100101101100000",
						 "101001111100101110010100",
						 "101001111100101111001000",
						 "101001111100101111111100",
						 "101001111100110000110000",
						 "101001111100110001100100",
						 "101001111100110010011000",
						 "101001111100100110001100",
						 "101001111100100110111111",
						 "101001111100100111110010",
						 "101001111100101000100101",
						 "101001111100101001011000",
						 "101001111100101010001011",
						 "101001111100101010111110",
						 "101001111100101011110001",
						 "101001111100101100100100",
						 "101001111100101101010111",
						 "101001111100101110001010",
						 "101001111100101110111101",
						 "101001111100101111110000",
						 "101001111100110000100011",
						 "101001111100110001010110",
						 "101001111100110010001001",
						 "101001111100100110001100",
						 "101001111100100110111111",
						 "101001111100100111110010",
						 "101001111100101000100101",
						 "101001111100101001011000",
						 "101001111100101010001011",
						 "101001111100101010111110",
						 "101001111100101011110001",
						 "101001111100101100100100",
						 "101001111100101101010111",
						 "101001111100101110001010",
						 "101001111100101110111101",
						 "101001111100101111110000",
						 "101001111100110000100011",
						 "101001111100110001010110",
						 "101001111100110010001001",
						 "101001111100100110001100",
						 "101001111100100110111111",
						 "101001111100100111110010",
						 "101001111100101000100101",
						 "101001111100101001011000",
						 "101001111100101010001011",
						 "101001111100101010111110",
						 "101001111100101011110001",
						 "101001111100101100100100",
						 "101001111100101101010111",
						 "101001111100101110001010",
						 "101001111100101110111101",
						 "101001111100101111110000",
						 "101001111100110000100011",
						 "101001111100110001010110",
						 "101001111100110010001001",
						 "101001111100100110001100",
						 "101001111100100110111110",
						 "101001111100100111110000",
						 "101001111100101000100010",
						 "101001111100101001010100",
						 "101001111100101010000110",
						 "101001111100101010111000",
						 "101001111100101011101010",
						 "101001111100101100011100",
						 "101001111100101101001110",
						 "101001111100101110000000",
						 "101001111100101110110010",
						 "101001111100101111100100",
						 "101001111100110000010110",
						 "101001111100110001001000",
						 "101001111100110001111010",
						 "101001111100100110001100",
						 "101001111100100110111110",
						 "101001111100100111110000",
						 "101001111100101000100010",
						 "101001111100101001010100",
						 "101001111100101010000110",
						 "101001111100101010111000",
						 "101001111100101011101010",
						 "101001111100101100011100",
						 "101001111100101101001110",
						 "101001111100101110000000",
						 "101001111100101110110010",
						 "101001111100101111100100",
						 "101001111100110000010110",
						 "101001111100110001001000",
						 "101001111100110001111010",
						 "101001111100100110001100",
						 "101001111100100110111110",
						 "101001111100100111110000",
						 "101001111100101000100010",
						 "101001111100101001010100",
						 "101001111100101010000110",
						 "101001111100101010111000",
						 "101001111100101011101010",
						 "101001111100101100011100",
						 "101001111100101101001110",
						 "101001111100101110000000",
						 "101001111100101110110010",
						 "101001111100101111100100",
						 "101001111100110000010110",
						 "101001111100110001001000",
						 "101001111100110001111010",
						 "101001111100100110001100",
						 "101001111100100110111101",
						 "101001111100100111101110",
						 "101001111100101000011111",
						 "101001111100101001010000",
						 "101001111100101010000001",
						 "101001111100101010110010",
						 "101001111100101011100011",
						 "101001111100101100010100",
						 "101001111100101101000101",
						 "101001111100101101110110",
						 "101001111100101110100111",
						 "101001111100101111011000",
						 "101001111100110000001001",
						 "101001111100110000111010",
						 "101001111100110001101011",
						 "101001111100100110001100",
						 "101001111100100110111101",
						 "101001111100100111101110",
						 "101001111100101000011111",
						 "101001111100101001010000",
						 "101001111100101010000001",
						 "101001111100101010110010",
						 "101001111100101011100011",
						 "101001111100101100010100",
						 "101001111100101101000101",
						 "101001111100101101110110",
						 "101001111100101110100111",
						 "101001111100101111011000",
						 "101001111100110000001001",
						 "101001111100110000111010",
						 "101001111100110001101011",
						 "101001111100100110001100",
						 "101001111100100110111100",
						 "101001111100100111101100",
						 "101001111100101000011100",
						 "101001111100101001001100",
						 "101001111100101001111100",
						 "101001111100101010101100",
						 "101001111100101011011100",
						 "101001111100101100001100",
						 "101001111100101100111100",
						 "101001111100101101101100",
						 "101001111100101110011100",
						 "101001111100101111001100",
						 "101001111100101111111100",
						 "101001111100110000101100",
						 "101001111100110001011100",
						 "101001111100100110001100",
						 "101001111100100110111100",
						 "101001111100100111101100",
						 "101001111100101000011100",
						 "101001111100101001001100",
						 "101001111100101001111100",
						 "101001111100101010101100",
						 "101001111100101011011100",
						 "101001111100101100001100",
						 "101001111100101100111100",
						 "101001111100101101101100",
						 "101001111100101110011100",
						 "101001111100101111001100",
						 "101001111100101111111100",
						 "101001111100110000101100",
						 "101001111100110001011100",
						 "101001111100100110001100",
						 "101001111100100110111100",
						 "101001111100100111101100",
						 "101001111100101000011100",
						 "101001111100101001001100",
						 "101001111100101001111100",
						 "101001111100101010101100",
						 "101001111100101011011100",
						 "101001111100101100001100",
						 "101001111100101100111100",
						 "101001111100101101101100",
						 "101001111100101110011100",
						 "101001111100101111001100",
						 "101001111100101111111100",
						 "101001111100110000101100",
						 "101001111100110001011100",
						 "101001111111001001001010",
						 "101001111111001001111001",
						 "101001111111001010101000",
						 "101001111111001011010111",
						 "101001111111001100000110",
						 "101001111111001100110101",
						 "101001111111001101100100",
						 "101001111111001110010011",
						 "101001111111001111000010",
						 "101001111111001111110001",
						 "101001111111010000100000",
						 "101001111111010001001111",
						 "101001111111010001111110",
						 "101001111111010010101101",
						 "101001111111010011011100",
						 "101001111111010100001011",
						 "101001111111001001001010",
						 "101001111111001001111001",
						 "101001111111001010101000",
						 "101001111111001011010111",
						 "101001111111001100000110",
						 "101001111111001100110101",
						 "101001111111001101100100",
						 "101001111111001110010011",
						 "101001111111001111000010",
						 "101001111111001111110001",
						 "101001111111010000100000",
						 "101001111111010001001111",
						 "101001111111010001111110",
						 "101001111111010010101101",
						 "101001111111010011011100",
						 "101001111111010100001011",
						 "101001111111001001001010",
						 "101001111111001001111000",
						 "101001111111001010100110",
						 "101001111111001011010100",
						 "101001111111001100000010",
						 "101001111111001100110000",
						 "101001111111001101011110",
						 "101001111111001110001100",
						 "101001111111001110111010",
						 "101001111111001111101000",
						 "101001111111010000010110",
						 "101001111111010001000100",
						 "101001111111010001110010",
						 "101001111111010010100000",
						 "101001111111010011001110",
						 "101001111111010011111100",
						 "101001111111001001001010",
						 "101001111111001001111000",
						 "101001111111001010100110",
						 "101001111111001011010100",
						 "101001111111001100000010",
						 "101001111111001100110000",
						 "101001111111001101011110",
						 "101001111111001110001100",
						 "101001111111001110111010",
						 "101001111111001111101000",
						 "101001111111010000010110",
						 "101001111111010001000100",
						 "101001111111010001110010",
						 "101001111111010010100000",
						 "101001111111010011001110",
						 "101001111111010011111100",
						 "101001111111001001001010",
						 "101001111111001001111000",
						 "101001111111001010100110",
						 "101001111111001011010100",
						 "101001111111001100000010",
						 "101001111111001100110000",
						 "101001111111001101011110",
						 "101001111111001110001100",
						 "101001111111001110111010",
						 "101001111111001111101000",
						 "101001111111010000010110",
						 "101001111111010001000100",
						 "101001111111010001110010",
						 "101001111111010010100000",
						 "101001111111010011001110",
						 "101001111111010011111100",
						 "101001111111001001001010",
						 "101001111111001001110111",
						 "101001111111001010100100",
						 "101001111111001011010001",
						 "101001111111001011111110",
						 "101001111111001100101011",
						 "101001111111001101011000",
						 "101001111111001110000101",
						 "101001111111001110110010",
						 "101001111111001111011111",
						 "101001111111010000001100",
						 "101001111111010000111001",
						 "101001111111010001100110",
						 "101001111111010010010011",
						 "101001111111010011000000",
						 "101001111111010011101101",
						 "101001111111001001001010",
						 "101001111111001001110111",
						 "101001111111001010100100",
						 "101001111111001011010001",
						 "101001111111001011111110",
						 "101001111111001100101011",
						 "101001111111001101011000",
						 "101001111111001110000101",
						 "101001111111001110110010",
						 "101001111111001111011111",
						 "101001111111010000001100",
						 "101001111111010000111001",
						 "101001111111010001100110",
						 "101001111111010010010011",
						 "101001111111010011000000",
						 "101001111111010011101101",
						 "101001111111001001001010",
						 "101001111111001001110111",
						 "101001111111001010100100",
						 "101001111111001011010001",
						 "101001111111001011111110",
						 "101001111111001100101011",
						 "101001111111001101011000",
						 "101001111111001110000101",
						 "101001111111001110110010",
						 "101001111111001111011111",
						 "101001111111010000001100",
						 "101001111111010000111001",
						 "101001111111010001100110",
						 "101001111111010010010011",
						 "101001111111010011000000",
						 "101001111111010011101101",
						 "101001111111001001001010",
						 "101001111111001001110110",
						 "101001111111001010100010",
						 "101001111111001011001110",
						 "101001111111001011111010",
						 "101001111111001100100110",
						 "101001111111001101010010",
						 "101001111111001101111110",
						 "101001111111001110101010",
						 "101001111111001111010110",
						 "101001111111010000000010",
						 "101001111111010000101110",
						 "101001111111010001011010",
						 "101001111111010010000110",
						 "101001111111010010110010",
						 "101001111111010011011110",
						 "101001111111001001001010",
						 "101001111111001001110110",
						 "101001111111001010100010",
						 "101001111111001011001110",
						 "101001111111001011111010",
						 "101001111111001100100110",
						 "101001111111001101010010",
						 "101001111111001101111110",
						 "101001111111001110101010",
						 "101001111111001111010110",
						 "101001111111010000000010",
						 "101001111111010000101110",
						 "101001111111010001011010",
						 "101001111111010010000110",
						 "101001111111010010110010",
						 "101001111111010011011110",
						 "101001111111001001001010",
						 "101001111111001001110101",
						 "101001111111001010100000",
						 "101001111111001011001011",
						 "101001111111001011110110",
						 "101001111111001100100001",
						 "101001111111001101001100",
						 "101001111111001101110111",
						 "101001111111001110100010",
						 "101001111111001111001101",
						 "101001111111001111111000",
						 "101001111111010000100011",
						 "101001111111010001001110",
						 "101001111111010001111001",
						 "101001111111010010100100",
						 "101001111111010011001111",
						 "101001111111001001001010",
						 "101001111111001001110101",
						 "101001111111001010100000",
						 "101001111111001011001011",
						 "101001111111001011110110",
						 "101001111111001100100001",
						 "101001111111001101001100",
						 "101001111111001101110111",
						 "101001111111001110100010",
						 "101001111111001111001101",
						 "101001111111001111111000",
						 "101001111111010000100011",
						 "101001111111010001001110",
						 "101001111111010001111001",
						 "101001111111010010100100",
						 "101001111111010011001111",
						 "101001111111001001001010",
						 "101001111111001001110101",
						 "101001111111001010100000",
						 "101001111111001011001011",
						 "101001111111001011110110",
						 "101001111111001100100001",
						 "101001111111001101001100",
						 "101001111111001101110111",
						 "101001111111001110100010",
						 "101001111111001111001101",
						 "101001111111001111111000",
						 "101001111111010000100011",
						 "101001111111010001001110",
						 "101001111111010001111001",
						 "101001111111010010100100",
						 "101001111111010011001111",
						 "101001111111001001001010",
						 "101001111111001001110100",
						 "101001111111001010011110",
						 "101001111111001011001000",
						 "101001111111001011110010",
						 "101001111111001100011100",
						 "101001111111001101000110",
						 "101001111111001101110000",
						 "101001111111001110011010",
						 "101001111111001111000100",
						 "101001111111001111101110",
						 "101001111111010000011000",
						 "101001111111010001000010",
						 "101001111111010001101100",
						 "101001111111010010010110",
						 "101001111111010011000000",
						 "101010000001101100001000",
						 "101010000001101100110010",
						 "101010000001101101011100",
						 "101010000001101110000110",
						 "101010000001101110110000",
						 "101010000001101111011010",
						 "101010000001110000000100",
						 "101010000001110000101110",
						 "101010000001110001011000",
						 "101010000001110010000010",
						 "101010000001110010101100",
						 "101010000001110011010110",
						 "101010000001110100000000",
						 "101010000001110100101010",
						 "101010000001110101010100",
						 "101010000001110101111110",
						 "101010000001101100001000",
						 "101010000001101100110001",
						 "101010000001101101011010",
						 "101010000001101110000011",
						 "101010000001101110101100",
						 "101010000001101111010101",
						 "101010000001101111111110",
						 "101010000001110000100111",
						 "101010000001110001010000",
						 "101010000001110001111001",
						 "101010000001110010100010",
						 "101010000001110011001011",
						 "101010000001110011110100",
						 "101010000001110100011101",
						 "101010000001110101000110",
						 "101010000001110101101111",
						 "101010000001101100001000",
						 "101010000001101100110001",
						 "101010000001101101011010",
						 "101010000001101110000011",
						 "101010000001101110101100",
						 "101010000001101111010101",
						 "101010000001101111111110",
						 "101010000001110000100111",
						 "101010000001110001010000",
						 "101010000001110001111001",
						 "101010000001110010100010",
						 "101010000001110011001011",
						 "101010000001110011110100",
						 "101010000001110100011101",
						 "101010000001110101000110",
						 "101010000001110101101111",
						 "101010000001101100001000",
						 "101010000001101100110001",
						 "101010000001101101011010",
						 "101010000001101110000011",
						 "101010000001101110101100",
						 "101010000001101111010101",
						 "101010000001101111111110",
						 "101010000001110000100111",
						 "101010000001110001010000",
						 "101010000001110001111001",
						 "101010000001110010100010",
						 "101010000001110011001011",
						 "101010000001110011110100",
						 "101010000001110100011101",
						 "101010000001110101000110",
						 "101010000001110101101111",
						 "101010000001101100001000",
						 "101010000001101100110000",
						 "101010000001101101011000",
						 "101010000001101110000000",
						 "101010000001101110101000",
						 "101010000001101111010000",
						 "101010000001101111111000",
						 "101010000001110000100000",
						 "101010000001110001001000",
						 "101010000001110001110000",
						 "101010000001110010011000",
						 "101010000001110011000000",
						 "101010000001110011101000",
						 "101010000001110100010000",
						 "101010000001110100111000",
						 "101010000001110101100000",
						 "101010000001101100001000",
						 "101010000001101100110000",
						 "101010000001101101011000",
						 "101010000001101110000000",
						 "101010000001101110101000",
						 "101010000001101111010000",
						 "101010000001101111111000",
						 "101010000001110000100000",
						 "101010000001110001001000",
						 "101010000001110001110000",
						 "101010000001110010011000",
						 "101010000001110011000000",
						 "101010000001110011101000",
						 "101010000001110100010000",
						 "101010000001110100111000",
						 "101010000001110101100000",
						 "101010000001101100001000",
						 "101010000001101100110000",
						 "101010000001101101011000",
						 "101010000001101110000000",
						 "101010000001101110101000",
						 "101010000001101111010000",
						 "101010000001101111111000",
						 "101010000001110000100000",
						 "101010000001110001001000",
						 "101010000001110001110000",
						 "101010000001110010011000",
						 "101010000001110011000000",
						 "101010000001110011101000",
						 "101010000001110100010000",
						 "101010000001110100111000",
						 "101010000001110101100000",
						 "101010000001101100001000",
						 "101010000001101100101111",
						 "101010000001101101010110",
						 "101010000001101101111101",
						 "101010000001101110100100",
						 "101010000001101111001011",
						 "101010000001101111110010",
						 "101010000001110000011001",
						 "101010000001110001000000",
						 "101010000001110001100111",
						 "101010000001110010001110",
						 "101010000001110010110101",
						 "101010000001110011011100",
						 "101010000001110100000011",
						 "101010000001110100101010",
						 "101010000001110101010001",
						 "101010000001101100001000",
						 "101010000001101100101111",
						 "101010000001101101010110",
						 "101010000001101101111101",
						 "101010000001101110100100",
						 "101010000001101111001011",
						 "101010000001101111110010",
						 "101010000001110000011001",
						 "101010000001110001000000",
						 "101010000001110001100111",
						 "101010000001110010001110",
						 "101010000001110010110101",
						 "101010000001110011011100",
						 "101010000001110100000011",
						 "101010000001110100101010",
						 "101010000001110101010001",
						 "101010000001101100001000",
						 "101010000001101100101110",
						 "101010000001101101010100",
						 "101010000001101101111010",
						 "101010000001101110100000",
						 "101010000001101111000110",
						 "101010000001101111101100",
						 "101010000001110000010010",
						 "101010000001110000111000",
						 "101010000001110001011110",
						 "101010000001110010000100",
						 "101010000001110010101010",
						 "101010000001110011010000",
						 "101010000001110011110110",
						 "101010000001110100011100",
						 "101010000001110101000010",
						 "101010000001101100001000",
						 "101010000001101100101110",
						 "101010000001101101010100",
						 "101010000001101101111010",
						 "101010000001101110100000",
						 "101010000001101111000110",
						 "101010000001101111101100",
						 "101010000001110000010010",
						 "101010000001110000111000",
						 "101010000001110001011110",
						 "101010000001110010000100",
						 "101010000001110010101010",
						 "101010000001110011010000",
						 "101010000001110011110110",
						 "101010000001110100011100",
						 "101010000001110101000010",
						 "101010000001101100001000",
						 "101010000001101100101110",
						 "101010000001101101010100",
						 "101010000001101101111010",
						 "101010000001101110100000",
						 "101010000001101111000110",
						 "101010000001101111101100",
						 "101010000001110000010010",
						 "101010000001110000111000",
						 "101010000001110001011110",
						 "101010000001110010000100",
						 "101010000001110010101010",
						 "101010000001110011010000",
						 "101010000001110011110110",
						 "101010000001110100011100",
						 "101010000001110101000010",
						 "101010000001101100001000",
						 "101010000001101100101101",
						 "101010000001101101010010",
						 "101010000001101101110111",
						 "101010000001101110011100",
						 "101010000001101111000001",
						 "101010000001101111100110",
						 "101010000001110000001011",
						 "101010000001110000110000",
						 "101010000001110001010101",
						 "101010000001110001111010",
						 "101010000001110010011111",
						 "101010000001110011000100",
						 "101010000001110011101001",
						 "101010000001110100001110",
						 "101010000001110100110011",
						 "101010000001101100001000",
						 "101010000001101100101101",
						 "101010000001101101010010",
						 "101010000001101101110111",
						 "101010000001101110011100",
						 "101010000001101111000001",
						 "101010000001101111100110",
						 "101010000001110000001011",
						 "101010000001110000110000",
						 "101010000001110001010101",
						 "101010000001110001111010",
						 "101010000001110010011111",
						 "101010000001110011000100",
						 "101010000001110011101001",
						 "101010000001110100001110",
						 "101010000001110100110011",
						 "101010000001101100001000",
						 "101010000001101100101100",
						 "101010000001101101010000",
						 "101010000001101101110100",
						 "101010000001101110011000",
						 "101010000001101110111100",
						 "101010000001101111100000",
						 "101010000001110000000100",
						 "101010000001110000101000",
						 "101010000001110001001100",
						 "101010000001110001110000",
						 "101010000001110010010100",
						 "101010000001110010111000",
						 "101010000001110011011100",
						 "101010000001110100000000",
						 "101010000001110100100100",
						 "101010000001101100001000",
						 "101010000001101100101100",
						 "101010000001101101010000",
						 "101010000001101101110100",
						 "101010000001101110011000",
						 "101010000001101110111100",
						 "101010000001101111100000",
						 "101010000001110000000100",
						 "101010000001110000101000",
						 "101010000001110001001100",
						 "101010000001110001110000",
						 "101010000001110010010100",
						 "101010000001110010111000",
						 "101010000001110011011100",
						 "101010000001110100000000",
						 "101010000001110100100100",
						 "101010000001101100001000",
						 "101010000001101100101100",
						 "101010000001101101010000",
						 "101010000001101101110100",
						 "101010000001101110011000",
						 "101010000001101110111100",
						 "101010000001101111100000",
						 "101010000001110000000100",
						 "101010000001110000101000",
						 "101010000001110001001100",
						 "101010000001110001110000",
						 "101010000001110010010100",
						 "101010000001110010111000",
						 "101010000001110011011100",
						 "101010000001110100000000",
						 "101010000001110100100100",
						 "101010000100001111000110",
						 "101010000100001111101001",
						 "101010000100010000001100",
						 "101010000100010000101111",
						 "101010000100010001010010",
						 "101010000100010001110101",
						 "101010000100010010011000",
						 "101010000100010010111011",
						 "101010000100010011011110",
						 "101010000100010100000001",
						 "101010000100010100100100",
						 "101010000100010101000111",
						 "101010000100010101101010",
						 "101010000100010110001101",
						 "101010000100010110110000",
						 "101010000100010111010011",
						 "101010000100001111000110",
						 "101010000100001111101001",
						 "101010000100010000001100",
						 "101010000100010000101111",
						 "101010000100010001010010",
						 "101010000100010001110101",
						 "101010000100010010011000",
						 "101010000100010010111011",
						 "101010000100010011011110",
						 "101010000100010100000001",
						 "101010000100010100100100",
						 "101010000100010101000111",
						 "101010000100010101101010",
						 "101010000100010110001101",
						 "101010000100010110110000",
						 "101010000100010111010011",
						 "101010000100001111000110",
						 "101010000100001111101001",
						 "101010000100010000001100",
						 "101010000100010000101111",
						 "101010000100010001010010",
						 "101010000100010001110101",
						 "101010000100010010011000",
						 "101010000100010010111011",
						 "101010000100010011011110",
						 "101010000100010100000001",
						 "101010000100010100100100",
						 "101010000100010101000111",
						 "101010000100010101101010",
						 "101010000100010110001101",
						 "101010000100010110110000",
						 "101010000100010111010011",
						 "101010000100001111000110",
						 "101010000100001111101000",
						 "101010000100010000001010",
						 "101010000100010000101100",
						 "101010000100010001001110",
						 "101010000100010001110000",
						 "101010000100010010010010",
						 "101010000100010010110100",
						 "101010000100010011010110",
						 "101010000100010011111000",
						 "101010000100010100011010",
						 "101010000100010100111100",
						 "101010000100010101011110",
						 "101010000100010110000000",
						 "101010000100010110100010",
						 "101010000100010111000100",
						 "101010000100001111000110",
						 "101010000100001111101000",
						 "101010000100010000001010",
						 "101010000100010000101100",
						 "101010000100010001001110",
						 "101010000100010001110000",
						 "101010000100010010010010",
						 "101010000100010010110100",
						 "101010000100010011010110",
						 "101010000100010011111000",
						 "101010000100010100011010",
						 "101010000100010100111100",
						 "101010000100010101011110",
						 "101010000100010110000000",
						 "101010000100010110100010",
						 "101010000100010111000100",
						 "101010000100001111000110",
						 "101010000100001111100111",
						 "101010000100010000001000",
						 "101010000100010000101001",
						 "101010000100010001001010",
						 "101010000100010001101011",
						 "101010000100010010001100",
						 "101010000100010010101101",
						 "101010000100010011001110",
						 "101010000100010011101111",
						 "101010000100010100010000",
						 "101010000100010100110001",
						 "101010000100010101010010",
						 "101010000100010101110011",
						 "101010000100010110010100",
						 "101010000100010110110101",
						 "101010000100001111000110",
						 "101010000100001111100111",
						 "101010000100010000001000",
						 "101010000100010000101001",
						 "101010000100010001001010",
						 "101010000100010001101011",
						 "101010000100010010001100",
						 "101010000100010010101101",
						 "101010000100010011001110",
						 "101010000100010011101111",
						 "101010000100010100010000",
						 "101010000100010100110001",
						 "101010000100010101010010",
						 "101010000100010101110011",
						 "101010000100010110010100",
						 "101010000100010110110101",
						 "101010000100001111000110",
						 "101010000100001111100111",
						 "101010000100010000001000",
						 "101010000100010000101001",
						 "101010000100010001001010",
						 "101010000100010001101011",
						 "101010000100010010001100",
						 "101010000100010010101101",
						 "101010000100010011001110",
						 "101010000100010011101111",
						 "101010000100010100010000",
						 "101010000100010100110001",
						 "101010000100010101010010",
						 "101010000100010101110011",
						 "101010000100010110010100",
						 "101010000100010110110101",
						 "101010000100001111000110",
						 "101010000100001111100110",
						 "101010000100010000000110",
						 "101010000100010000100110",
						 "101010000100010001000110",
						 "101010000100010001100110",
						 "101010000100010010000110",
						 "101010000100010010100110",
						 "101010000100010011000110",
						 "101010000100010011100110",
						 "101010000100010100000110",
						 "101010000100010100100110",
						 "101010000100010101000110",
						 "101010000100010101100110",
						 "101010000100010110000110",
						 "101010000100010110100110",
						 "101010000100001111000110",
						 "101010000100001111100110",
						 "101010000100010000000110",
						 "101010000100010000100110",
						 "101010000100010001000110",
						 "101010000100010001100110",
						 "101010000100010010000110",
						 "101010000100010010100110",
						 "101010000100010011000110",
						 "101010000100010011100110",
						 "101010000100010100000110",
						 "101010000100010100100110",
						 "101010000100010101000110",
						 "101010000100010101100110",
						 "101010000100010110000110",
						 "101010000100010110100110",
						 "101010000100001111000110",
						 "101010000100001111100101",
						 "101010000100010000000100",
						 "101010000100010000100011",
						 "101010000100010001000010",
						 "101010000100010001100001",
						 "101010000100010010000000",
						 "101010000100010010011111",
						 "101010000100010010111110",
						 "101010000100010011011101",
						 "101010000100010011111100",
						 "101010000100010100011011",
						 "101010000100010100111010",
						 "101010000100010101011001",
						 "101010000100010101111000",
						 "101010000100010110010111",
						 "101010000100001111000110",
						 "101010000100001111100101",
						 "101010000100010000000100",
						 "101010000100010000100011",
						 "101010000100010001000010",
						 "101010000100010001100001",
						 "101010000100010010000000",
						 "101010000100010010011111",
						 "101010000100010010111110",
						 "101010000100010011011101",
						 "101010000100010011111100",
						 "101010000100010100011011",
						 "101010000100010100111010",
						 "101010000100010101011001",
						 "101010000100010101111000",
						 "101010000100010110010111",
						 "101010000100001111000110",
						 "101010000100001111100101",
						 "101010000100010000000100",
						 "101010000100010000100011",
						 "101010000100010001000010",
						 "101010000100010001100001",
						 "101010000100010010000000",
						 "101010000100010010011111",
						 "101010000100010010111110",
						 "101010000100010011011101",
						 "101010000100010011111100",
						 "101010000100010100011011",
						 "101010000100010100111010",
						 "101010000100010101011001",
						 "101010000100010101111000",
						 "101010000100010110010111",
						 "101010000100001111000110",
						 "101010000100001111100100",
						 "101010000100010000000010",
						 "101010000100010000100000",
						 "101010000100010000111110",
						 "101010000100010001011100",
						 "101010000100010001111010",
						 "101010000100010010011000",
						 "101010000100010010110110",
						 "101010000100010011010100",
						 "101010000100010011110010",
						 "101010000100010100010000",
						 "101010000100010100101110",
						 "101010000100010101001100",
						 "101010000100010101101010",
						 "101010000100010110001000",
						 "101010000100001111000110",
						 "101010000100001111100100",
						 "101010000100010000000010",
						 "101010000100010000100000",
						 "101010000100010000111110",
						 "101010000100010001011100",
						 "101010000100010001111010",
						 "101010000100010010011000",
						 "101010000100010010110110",
						 "101010000100010011010100",
						 "101010000100010011110010",
						 "101010000100010100010000",
						 "101010000100010100101110",
						 "101010000100010101001100",
						 "101010000100010101101010",
						 "101010000100010110001000",
						 "101010000100001111000110",
						 "101010000100001111100011",
						 "101010000100010000000000",
						 "101010000100010000011101",
						 "101010000100010000111010",
						 "101010000100010001010111",
						 "101010000100010001110100",
						 "101010000100010010010001",
						 "101010000100010010101110",
						 "101010000100010011001011",
						 "101010000100010011101000",
						 "101010000100010100000101",
						 "101010000100010100100010",
						 "101010000100010100111111",
						 "101010000100010101011100",
						 "101010000100010101111001",
						 "101010000100001111000110",
						 "101010000100001111100011",
						 "101010000100010000000000",
						 "101010000100010000011101",
						 "101010000100010000111010",
						 "101010000100010001010111",
						 "101010000100010001110100",
						 "101010000100010010010001",
						 "101010000100010010101110",
						 "101010000100010011001011",
						 "101010000100010011101000",
						 "101010000100010100000101",
						 "101010000100010100100010",
						 "101010000100010100111111",
						 "101010000100010101011100",
						 "101010000100010101111001",
						 "101010000100001111000110",
						 "101010000100001111100011",
						 "101010000100010000000000",
						 "101010000100010000011101",
						 "101010000100010000111010",
						 "101010000100010001010111",
						 "101010000100010001110100",
						 "101010000100010010010001",
						 "101010000100010010101110",
						 "101010000100010011001011",
						 "101010000100010011101000",
						 "101010000100010100000101",
						 "101010000100010100100010",
						 "101010000100010100111111",
						 "101010000100010101011100",
						 "101010000100010101111001",
						 "101010000100001111000110",
						 "101010000100001111100010",
						 "101010000100001111111110",
						 "101010000100010000011010",
						 "101010000100010000110110",
						 "101010000100010001010010",
						 "101010000100010001101110",
						 "101010000100010010001010",
						 "101010000100010010100110",
						 "101010000100010011000010",
						 "101010000100010011011110",
						 "101010000100010011111010",
						 "101010000100010100010110",
						 "101010000100010100110010",
						 "101010000100010101001110",
						 "101010000100010101101010",
						 "101010000100001111000110",
						 "101010000100001111100010",
						 "101010000100001111111110",
						 "101010000100010000011010",
						 "101010000100010000110110",
						 "101010000100010001010010",
						 "101010000100010001101110",
						 "101010000100010010001010",
						 "101010000100010010100110",
						 "101010000100010011000010",
						 "101010000100010011011110",
						 "101010000100010011111010",
						 "101010000100010100010110",
						 "101010000100010100110010",
						 "101010000100010101001110",
						 "101010000100010101101010",
						 "101010000100001111000110",
						 "101010000100001111100010",
						 "101010000100001111111110",
						 "101010000100010000011010",
						 "101010000100010000110110",
						 "101010000100010001010010",
						 "101010000100010001101110",
						 "101010000100010010001010",
						 "101010000100010010100110",
						 "101010000100010011000010",
						 "101010000100010011011110",
						 "101010000100010011111010",
						 "101010000100010100010110",
						 "101010000100010100110010",
						 "101010000100010101001110",
						 "101010000100010101101010",
						 "101010000110110010000100",
						 "101010000110110010011111",
						 "101010000110110010111010",
						 "101010000110110011010101",
						 "101010000110110011110000",
						 "101010000110110100001011",
						 "101010000110110100100110",
						 "101010000110110101000001",
						 "101010000110110101011100",
						 "101010000110110101110111",
						 "101010000110110110010010",
						 "101010000110110110101101",
						 "101010000110110111001000",
						 "101010000110110111100011",
						 "101010000110110111111110",
						 "101010000110111000011001",
						 "101010000110110010000100",
						 "101010000110110010011111",
						 "101010000110110010111010",
						 "101010000110110011010101",
						 "101010000110110011110000",
						 "101010000110110100001011",
						 "101010000110110100100110",
						 "101010000110110101000001",
						 "101010000110110101011100",
						 "101010000110110101110111",
						 "101010000110110110010010",
						 "101010000110110110101101",
						 "101010000110110111001000",
						 "101010000110110111100011",
						 "101010000110110111111110",
						 "101010000110111000011001",
						 "101010000110110010000100",
						 "101010000110110010011110",
						 "101010000110110010111000",
						 "101010000110110011010010",
						 "101010000110110011101100",
						 "101010000110110100000110",
						 "101010000110110100100000",
						 "101010000110110100111010",
						 "101010000110110101010100",
						 "101010000110110101101110",
						 "101010000110110110001000",
						 "101010000110110110100010",
						 "101010000110110110111100",
						 "101010000110110111010110",
						 "101010000110110111110000",
						 "101010000110111000001010",
						 "101010000110110010000100",
						 "101010000110110010011110",
						 "101010000110110010111000",
						 "101010000110110011010010",
						 "101010000110110011101100",
						 "101010000110110100000110",
						 "101010000110110100100000",
						 "101010000110110100111010",
						 "101010000110110101010100",
						 "101010000110110101101110",
						 "101010000110110110001000",
						 "101010000110110110100010",
						 "101010000110110110111100",
						 "101010000110110111010110",
						 "101010000110110111110000",
						 "101010000110111000001010",
						 "101010000110110010000100",
						 "101010000110110010011110",
						 "101010000110110010111000",
						 "101010000110110011010010",
						 "101010000110110011101100",
						 "101010000110110100000110",
						 "101010000110110100100000",
						 "101010000110110100111010",
						 "101010000110110101010100",
						 "101010000110110101101110",
						 "101010000110110110001000",
						 "101010000110110110100010",
						 "101010000110110110111100",
						 "101010000110110111010110",
						 "101010000110110111110000",
						 "101010000110111000001010",
						 "101010000110110010000100",
						 "101010000110110010011101",
						 "101010000110110010110110",
						 "101010000110110011001111",
						 "101010000110110011101000",
						 "101010000110110100000001",
						 "101010000110110100011010",
						 "101010000110110100110011",
						 "101010000110110101001100",
						 "101010000110110101100101",
						 "101010000110110101111110",
						 "101010000110110110010111",
						 "101010000110110110110000",
						 "101010000110110111001001",
						 "101010000110110111100010",
						 "101010000110110111111011",
						 "101010000110110010000100",
						 "101010000110110010011101",
						 "101010000110110010110110",
						 "101010000110110011001111",
						 "101010000110110011101000",
						 "101010000110110100000001",
						 "101010000110110100011010",
						 "101010000110110100110011",
						 "101010000110110101001100",
						 "101010000110110101100101",
						 "101010000110110101111110",
						 "101010000110110110010111",
						 "101010000110110110110000",
						 "101010000110110111001001",
						 "101010000110110111100010",
						 "101010000110110111111011",
						 "101010000110110010000100",
						 "101010000110110010011100",
						 "101010000110110010110100",
						 "101010000110110011001100",
						 "101010000110110011100100",
						 "101010000110110011111100",
						 "101010000110110100010100",
						 "101010000110110100101100",
						 "101010000110110101000100",
						 "101010000110110101011100",
						 "101010000110110101110100",
						 "101010000110110110001100",
						 "101010000110110110100100",
						 "101010000110110110111100",
						 "101010000110110111010100",
						 "101010000110110111101100",
						 "101010000110110010000100",
						 "101010000110110010011100",
						 "101010000110110010110100",
						 "101010000110110011001100",
						 "101010000110110011100100",
						 "101010000110110011111100",
						 "101010000110110100010100",
						 "101010000110110100101100",
						 "101010000110110101000100",
						 "101010000110110101011100",
						 "101010000110110101110100",
						 "101010000110110110001100",
						 "101010000110110110100100",
						 "101010000110110110111100",
						 "101010000110110111010100",
						 "101010000110110111101100",
						 "101010000110110010000100",
						 "101010000110110010011100",
						 "101010000110110010110100",
						 "101010000110110011001100",
						 "101010000110110011100100",
						 "101010000110110011111100",
						 "101010000110110100010100",
						 "101010000110110100101100",
						 "101010000110110101000100",
						 "101010000110110101011100",
						 "101010000110110101110100",
						 "101010000110110110001100",
						 "101010000110110110100100",
						 "101010000110110110111100",
						 "101010000110110111010100",
						 "101010000110110111101100",
						 "101010000110110010000100",
						 "101010000110110010011011",
						 "101010000110110010110010",
						 "101010000110110011001001",
						 "101010000110110011100000",
						 "101010000110110011110111",
						 "101010000110110100001110",
						 "101010000110110100100101",
						 "101010000110110100111100",
						 "101010000110110101010011",
						 "101010000110110101101010",
						 "101010000110110110000001",
						 "101010000110110110011000",
						 "101010000110110110101111",
						 "101010000110110111000110",
						 "101010000110110111011101",
						 "101010000110110010000100",
						 "101010000110110010011011",
						 "101010000110110010110010",
						 "101010000110110011001001",
						 "101010000110110011100000",
						 "101010000110110011110111",
						 "101010000110110100001110",
						 "101010000110110100100101",
						 "101010000110110100111100",
						 "101010000110110101010011",
						 "101010000110110101101010",
						 "101010000110110110000001",
						 "101010000110110110011000",
						 "101010000110110110101111",
						 "101010000110110111000110",
						 "101010000110110111011101",
						 "101010000110110010000100",
						 "101010000110110010011010",
						 "101010000110110010110000",
						 "101010000110110011000110",
						 "101010000110110011011100",
						 "101010000110110011110010",
						 "101010000110110100001000",
						 "101010000110110100011110",
						 "101010000110110100110100",
						 "101010000110110101001010",
						 "101010000110110101100000",
						 "101010000110110101110110",
						 "101010000110110110001100",
						 "101010000110110110100010",
						 "101010000110110110111000",
						 "101010000110110111001110",
						 "101010000110110010000100",
						 "101010000110110010011010",
						 "101010000110110010110000",
						 "101010000110110011000110",
						 "101010000110110011011100",
						 "101010000110110011110010",
						 "101010000110110100001000",
						 "101010000110110100011110",
						 "101010000110110100110100",
						 "101010000110110101001010",
						 "101010000110110101100000",
						 "101010000110110101110110",
						 "101010000110110110001100",
						 "101010000110110110100010",
						 "101010000110110110111000",
						 "101010000110110111001110",
						 "101010000110110010000100",
						 "101010000110110010011010",
						 "101010000110110010110000",
						 "101010000110110011000110",
						 "101010000110110011011100",
						 "101010000110110011110010",
						 "101010000110110100001000",
						 "101010000110110100011110",
						 "101010000110110100110100",
						 "101010000110110101001010",
						 "101010000110110101100000",
						 "101010000110110101110110",
						 "101010000110110110001100",
						 "101010000110110110100010",
						 "101010000110110110111000",
						 "101010000110110111001110",
						 "101010000110110010000100",
						 "101010000110110010011001",
						 "101010000110110010101110",
						 "101010000110110011000011",
						 "101010000110110011011000",
						 "101010000110110011101101",
						 "101010000110110100000010",
						 "101010000110110100010111",
						 "101010000110110100101100",
						 "101010000110110101000001",
						 "101010000110110101010110",
						 "101010000110110101101011",
						 "101010000110110110000000",
						 "101010000110110110010101",
						 "101010000110110110101010",
						 "101010000110110110111111",
						 "101010000110110010000100",
						 "101010000110110010011001",
						 "101010000110110010101110",
						 "101010000110110011000011",
						 "101010000110110011011000",
						 "101010000110110011101101",
						 "101010000110110100000010",
						 "101010000110110100010111",
						 "101010000110110100101100",
						 "101010000110110101000001",
						 "101010000110110101010110",
						 "101010000110110101101011",
						 "101010000110110110000000",
						 "101010000110110110010101",
						 "101010000110110110101010",
						 "101010000110110110111111",
						 "101010000110110010000100",
						 "101010000110110010011001",
						 "101010000110110010101110",
						 "101010000110110011000011",
						 "101010000110110011011000",
						 "101010000110110011101101",
						 "101010000110110100000010",
						 "101010000110110100010111",
						 "101010000110110100101100",
						 "101010000110110101000001",
						 "101010000110110101010110",
						 "101010000110110101101011",
						 "101010000110110110000000",
						 "101010000110110110010101",
						 "101010000110110110101010",
						 "101010000110110110111111",
						 "101010000110110010000100",
						 "101010000110110010011000",
						 "101010000110110010101100",
						 "101010000110110011000000",
						 "101010000110110011010100",
						 "101010000110110011101000",
						 "101010000110110011111100",
						 "101010000110110100010000",
						 "101010000110110100100100",
						 "101010000110110100111000",
						 "101010000110110101001100",
						 "101010000110110101100000",
						 "101010000110110101110100",
						 "101010000110110110001000",
						 "101010000110110110011100",
						 "101010000110110110110000",
						 "101010000110110010000100",
						 "101010000110110010011000",
						 "101010000110110010101100",
						 "101010000110110011000000",
						 "101010000110110011010100",
						 "101010000110110011101000",
						 "101010000110110011111100",
						 "101010000110110100010000",
						 "101010000110110100100100",
						 "101010000110110100111000",
						 "101010000110110101001100",
						 "101010000110110101100000",
						 "101010000110110101110100",
						 "101010000110110110001000",
						 "101010000110110110011100",
						 "101010000110110110110000",
						 "101010000110110010000100",
						 "101010000110110010010111",
						 "101010000110110010101010",
						 "101010000110110010111101",
						 "101010000110110011010000",
						 "101010000110110011100011",
						 "101010000110110011110110",
						 "101010000110110100001001",
						 "101010000110110100011100",
						 "101010000110110100101111",
						 "101010000110110101000010",
						 "101010000110110101010101",
						 "101010000110110101101000",
						 "101010000110110101111011",
						 "101010000110110110001110",
						 "101010000110110110100001",
						 "101010000110110010000100",
						 "101010000110110010010111",
						 "101010000110110010101010",
						 "101010000110110010111101",
						 "101010000110110011010000",
						 "101010000110110011100011",
						 "101010000110110011110110",
						 "101010000110110100001001",
						 "101010000110110100011100",
						 "101010000110110100101111",
						 "101010000110110101000010",
						 "101010000110110101010101",
						 "101010000110110101101000",
						 "101010000110110101111011",
						 "101010000110110110001110",
						 "101010000110110110100001",
						 "101010000110110010000100",
						 "101010000110110010010111",
						 "101010000110110010101010",
						 "101010000110110010111101",
						 "101010000110110011010000",
						 "101010000110110011100011",
						 "101010000110110011110110",
						 "101010000110110100001001",
						 "101010000110110100011100",
						 "101010000110110100101111",
						 "101010000110110101000010",
						 "101010000110110101010101",
						 "101010000110110101101000",
						 "101010000110110101111011",
						 "101010000110110110001110",
						 "101010000110110110100001",
						 "101010000110110010000100",
						 "101010000110110010010110",
						 "101010000110110010101000",
						 "101010000110110010111010",
						 "101010000110110011001100",
						 "101010000110110011011110",
						 "101010000110110011110000",
						 "101010000110110100000010",
						 "101010000110110100010100",
						 "101010000110110100100110",
						 "101010000110110100111000",
						 "101010000110110101001010",
						 "101010000110110101011100",
						 "101010000110110101101110",
						 "101010000110110110000000",
						 "101010000110110110010010",
						 "101010000110110010000100",
						 "101010000110110010010110",
						 "101010000110110010101000",
						 "101010000110110010111010",
						 "101010000110110011001100",
						 "101010000110110011011110",
						 "101010000110110011110000",
						 "101010000110110100000010",
						 "101010000110110100010100",
						 "101010000110110100100110",
						 "101010000110110100111000",
						 "101010000110110101001010",
						 "101010000110110101011100",
						 "101010000110110101101110",
						 "101010000110110110000000",
						 "101010000110110110010010",
						 "101010000110110010000100",
						 "101010000110110010010101",
						 "101010000110110010100110",
						 "101010000110110010110111",
						 "101010000110110011001000",
						 "101010000110110011011001",
						 "101010000110110011101010",
						 "101010000110110011111011",
						 "101010000110110100001100",
						 "101010000110110100011101",
						 "101010000110110100101110",
						 "101010000110110100111111",
						 "101010000110110101010000",
						 "101010000110110101100001",
						 "101010000110110101110010",
						 "101010000110110110000011",
						 "101010000110110010000100",
						 "101010000110110010010101",
						 "101010000110110010100110",
						 "101010000110110010110111",
						 "101010000110110011001000",
						 "101010000110110011011001",
						 "101010000110110011101010",
						 "101010000110110011111011",
						 "101010000110110100001100",
						 "101010000110110100011101",
						 "101010000110110100101110",
						 "101010000110110100111111",
						 "101010000110110101010000",
						 "101010000110110101100001",
						 "101010000110110101110010",
						 "101010000110110110000011",
						 "101010000110110010000100",
						 "101010000110110010010101",
						 "101010000110110010100110",
						 "101010000110110010110111",
						 "101010000110110011001000",
						 "101010000110110011011001",
						 "101010000110110011101010",
						 "101010000110110011111011",
						 "101010000110110100001100",
						 "101010000110110100011101",
						 "101010000110110100101110",
						 "101010000110110100111111",
						 "101010000110110101010000",
						 "101010000110110101100001",
						 "101010000110110101110010",
						 "101010000110110110000011",
						 "101010000110110010000100",
						 "101010000110110010010100",
						 "101010000110110010100100",
						 "101010000110110010110100",
						 "101010000110110011000100",
						 "101010000110110011010100",
						 "101010000110110011100100",
						 "101010000110110011110100",
						 "101010000110110100000100",
						 "101010000110110100010100",
						 "101010000110110100100100",
						 "101010000110110100110100",
						 "101010000110110101000100",
						 "101010000110110101010100",
						 "101010000110110101100100",
						 "101010000110110101110100",
						 "101010000110110010000100",
						 "101010000110110010010100",
						 "101010000110110010100100",
						 "101010000110110010110100",
						 "101010000110110011000100",
						 "101010000110110011010100",
						 "101010000110110011100100",
						 "101010000110110011110100",
						 "101010000110110100000100",
						 "101010000110110100010100",
						 "101010000110110100100100",
						 "101010000110110100110100",
						 "101010000110110101000100",
						 "101010000110110101010100",
						 "101010000110110101100100",
						 "101010000110110101110100",
						 "101010001001010101000010",
						 "101010001001010101010001",
						 "101010001001010101100000",
						 "101010001001010101101111",
						 "101010001001010101111110",
						 "101010001001010110001101",
						 "101010001001010110011100",
						 "101010001001010110101011",
						 "101010001001010110111010",
						 "101010001001010111001001",
						 "101010001001010111011000",
						 "101010001001010111100111",
						 "101010001001010111110110",
						 "101010001001011000000101",
						 "101010001001011000010100",
						 "101010001001011000100011",
						 "101010001001010101000010",
						 "101010001001010101010001",
						 "101010001001010101100000",
						 "101010001001010101101111",
						 "101010001001010101111110",
						 "101010001001010110001101",
						 "101010001001010110011100",
						 "101010001001010110101011",
						 "101010001001010110111010",
						 "101010001001010111001001",
						 "101010001001010111011000",
						 "101010001001010111100111",
						 "101010001001010111110110",
						 "101010001001011000000101",
						 "101010001001011000010100",
						 "101010001001011000100011",
						 "101010001001010101000010",
						 "101010001001010101010001",
						 "101010001001010101100000",
						 "101010001001010101101111",
						 "101010001001010101111110",
						 "101010001001010110001101",
						 "101010001001010110011100",
						 "101010001001010110101011",
						 "101010001001010110111010",
						 "101010001001010111001001",
						 "101010001001010111011000",
						 "101010001001010111100111",
						 "101010001001010111110110",
						 "101010001001011000000101",
						 "101010001001011000010100",
						 "101010001001011000100011",
						 "101010001001010101000010",
						 "101010001001010101010000",
						 "101010001001010101011110",
						 "101010001001010101101100",
						 "101010001001010101111010",
						 "101010001001010110001000",
						 "101010001001010110010110",
						 "101010001001010110100100",
						 "101010001001010110110010",
						 "101010001001010111000000",
						 "101010001001010111001110",
						 "101010001001010111011100",
						 "101010001001010111101010",
						 "101010001001010111111000",
						 "101010001001011000000110",
						 "101010001001011000010100",
						 "101010001001010101000010",
						 "101010001001010101010000",
						 "101010001001010101011110",
						 "101010001001010101101100",
						 "101010001001010101111010",
						 "101010001001010110001000",
						 "101010001001010110010110",
						 "101010001001010110100100",
						 "101010001001010110110010",
						 "101010001001010111000000",
						 "101010001001010111001110",
						 "101010001001010111011100",
						 "101010001001010111101010",
						 "101010001001010111111000",
						 "101010001001011000000110",
						 "101010001001011000010100",
						 "101010001001010101000010",
						 "101010001001010101001111",
						 "101010001001010101011100",
						 "101010001001010101101001",
						 "101010001001010101110110",
						 "101010001001010110000011",
						 "101010001001010110010000",
						 "101010001001010110011101",
						 "101010001001010110101010",
						 "101010001001010110110111",
						 "101010001001010111000100",
						 "101010001001010111010001",
						 "101010001001010111011110",
						 "101010001001010111101011",
						 "101010001001010111111000",
						 "101010001001011000000101",
						 "101010001001010101000010",
						 "101010001001010101001111",
						 "101010001001010101011100",
						 "101010001001010101101001",
						 "101010001001010101110110",
						 "101010001001010110000011",
						 "101010001001010110010000",
						 "101010001001010110011101",
						 "101010001001010110101010",
						 "101010001001010110110111",
						 "101010001001010111000100",
						 "101010001001010111010001",
						 "101010001001010111011110",
						 "101010001001010111101011",
						 "101010001001010111111000",
						 "101010001001011000000101",
						 "101010001001010101000010",
						 "101010001001010101001111",
						 "101010001001010101011100",
						 "101010001001010101101001",
						 "101010001001010101110110",
						 "101010001001010110000011",
						 "101010001001010110010000",
						 "101010001001010110011101",
						 "101010001001010110101010",
						 "101010001001010110110111",
						 "101010001001010111000100",
						 "101010001001010111010001",
						 "101010001001010111011110",
						 "101010001001010111101011",
						 "101010001001010111111000",
						 "101010001001011000000101",
						 "101010001001010101000010",
						 "101010001001010101001110",
						 "101010001001010101011010",
						 "101010001001010101100110",
						 "101010001001010101110010",
						 "101010001001010101111110",
						 "101010001001010110001010",
						 "101010001001010110010110",
						 "101010001001010110100010",
						 "101010001001010110101110",
						 "101010001001010110111010",
						 "101010001001010111000110",
						 "101010001001010111010010",
						 "101010001001010111011110",
						 "101010001001010111101010",
						 "101010001001010111110110",
						 "101010001001010101000010",
						 "101010001001010101001110",
						 "101010001001010101011010",
						 "101010001001010101100110",
						 "101010001001010101110010",
						 "101010001001010101111110",
						 "101010001001010110001010",
						 "101010001001010110010110",
						 "101010001001010110100010",
						 "101010001001010110101110",
						 "101010001001010110111010",
						 "101010001001010111000110",
						 "101010001001010111010010",
						 "101010001001010111011110",
						 "101010001001010111101010",
						 "101010001001010111110110",
						 "101010001001010101000010",
						 "101010001001010101001110",
						 "101010001001010101011010",
						 "101010001001010101100110",
						 "101010001001010101110010",
						 "101010001001010101111110",
						 "101010001001010110001010",
						 "101010001001010110010110",
						 "101010001001010110100010",
						 "101010001001010110101110",
						 "101010001001010110111010",
						 "101010001001010111000110",
						 "101010001001010111010010",
						 "101010001001010111011110",
						 "101010001001010111101010",
						 "101010001001010111110110",
						 "101010001001010101000010",
						 "101010001001010101001101",
						 "101010001001010101011000",
						 "101010001001010101100011",
						 "101010001001010101101110",
						 "101010001001010101111001",
						 "101010001001010110000100",
						 "101010001001010110001111",
						 "101010001001010110011010",
						 "101010001001010110100101",
						 "101010001001010110110000",
						 "101010001001010110111011",
						 "101010001001010111000110",
						 "101010001001010111010001",
						 "101010001001010111011100",
						 "101010001001010111100111",
						 "101010001001010101000010",
						 "101010001001010101001101",
						 "101010001001010101011000",
						 "101010001001010101100011",
						 "101010001001010101101110",
						 "101010001001010101111001",
						 "101010001001010110000100",
						 "101010001001010110001111",
						 "101010001001010110011010",
						 "101010001001010110100101",
						 "101010001001010110110000",
						 "101010001001010110111011",
						 "101010001001010111000110",
						 "101010001001010111010001",
						 "101010001001010111011100",
						 "101010001001010111100111",
						 "101010001001010101000010",
						 "101010001001010101001100",
						 "101010001001010101010110",
						 "101010001001010101100000",
						 "101010001001010101101010",
						 "101010001001010101110100",
						 "101010001001010101111110",
						 "101010001001010110001000",
						 "101010001001010110010010",
						 "101010001001010110011100",
						 "101010001001010110100110",
						 "101010001001010110110000",
						 "101010001001010110111010",
						 "101010001001010111000100",
						 "101010001001010111001110",
						 "101010001001010111011000",
						 "101010001001010101000010",
						 "101010001001010101001100",
						 "101010001001010101010110",
						 "101010001001010101100000",
						 "101010001001010101101010",
						 "101010001001010101110100",
						 "101010001001010101111110",
						 "101010001001010110001000",
						 "101010001001010110010010",
						 "101010001001010110011100",
						 "101010001001010110100110",
						 "101010001001010110110000",
						 "101010001001010110111010",
						 "101010001001010111000100",
						 "101010001001010111001110",
						 "101010001001010111011000",
						 "101010001001010101000010",
						 "101010001001010101001100",
						 "101010001001010101010110",
						 "101010001001010101100000",
						 "101010001001010101101010",
						 "101010001001010101110100",
						 "101010001001010101111110",
						 "101010001001010110001000",
						 "101010001001010110010010",
						 "101010001001010110011100",
						 "101010001001010110100110",
						 "101010001001010110110000",
						 "101010001001010110111010",
						 "101010001001010111000100",
						 "101010001001010111001110",
						 "101010001001010111011000",
						 "101010001001010101000010",
						 "101010001001010101001011",
						 "101010001001010101010100",
						 "101010001001010101011101",
						 "101010001001010101100110",
						 "101010001001010101101111",
						 "101010001001010101111000",
						 "101010001001010110000001",
						 "101010001001010110001010",
						 "101010001001010110010011",
						 "101010001001010110011100",
						 "101010001001010110100101",
						 "101010001001010110101110",
						 "101010001001010110110111",
						 "101010001001010111000000",
						 "101010001001010111001001",
						 "101010001001010101000010",
						 "101010001001010101001011",
						 "101010001001010101010100",
						 "101010001001010101011101",
						 "101010001001010101100110",
						 "101010001001010101101111",
						 "101010001001010101111000",
						 "101010001001010110000001",
						 "101010001001010110001010",
						 "101010001001010110010011",
						 "101010001001010110011100",
						 "101010001001010110100101",
						 "101010001001010110101110",
						 "101010001001010110110111",
						 "101010001001010111000000",
						 "101010001001010111001001",
						 "101010001001010101000010",
						 "101010001001010101001010",
						 "101010001001010101010010",
						 "101010001001010101011010",
						 "101010001001010101100010",
						 "101010001001010101101010",
						 "101010001001010101110010",
						 "101010001001010101111010",
						 "101010001001010110000010",
						 "101010001001010110001010",
						 "101010001001010110010010",
						 "101010001001010110011010",
						 "101010001001010110100010",
						 "101010001001010110101010",
						 "101010001001010110110010",
						 "101010001001010110111010",
						 "101010001001010101000010",
						 "101010001001010101001010",
						 "101010001001010101010010",
						 "101010001001010101011010",
						 "101010001001010101100010",
						 "101010001001010101101010",
						 "101010001001010101110010",
						 "101010001001010101111010",
						 "101010001001010110000010",
						 "101010001001010110001010",
						 "101010001001010110010010",
						 "101010001001010110011010",
						 "101010001001010110100010",
						 "101010001001010110101010",
						 "101010001001010110110010",
						 "101010001001010110111010",
						 "101010001001010101000010",
						 "101010001001010101001010",
						 "101010001001010101010010",
						 "101010001001010101011010",
						 "101010001001010101100010",
						 "101010001001010101101010",
						 "101010001001010101110010",
						 "101010001001010101111010",
						 "101010001001010110000010",
						 "101010001001010110001010",
						 "101010001001010110010010",
						 "101010001001010110011010",
						 "101010001001010110100010",
						 "101010001001010110101010",
						 "101010001001010110110010",
						 "101010001001010110111010",
						 "101010001001010101000010",
						 "101010001001010101001001",
						 "101010001001010101010000",
						 "101010001001010101010111",
						 "101010001001010101011110",
						 "101010001001010101100101",
						 "101010001001010101101100",
						 "101010001001010101110011",
						 "101010001001010101111010",
						 "101010001001010110000001",
						 "101010001001010110001000",
						 "101010001001010110001111",
						 "101010001001010110010110",
						 "101010001001010110011101",
						 "101010001001010110100100",
						 "101010001001010110101011",
						 "101010001001010101000010",
						 "101010001001010101001001",
						 "101010001001010101010000",
						 "101010001001010101010111",
						 "101010001001010101011110",
						 "101010001001010101100101",
						 "101010001001010101101100",
						 "101010001001010101110011",
						 "101010001001010101111010",
						 "101010001001010110000001",
						 "101010001001010110001000",
						 "101010001001010110001111",
						 "101010001001010110010110",
						 "101010001001010110011101",
						 "101010001001010110100100",
						 "101010001001010110101011",
						 "101010001001010101000010",
						 "101010001001010101001000",
						 "101010001001010101001110",
						 "101010001001010101010100",
						 "101010001001010101011010",
						 "101010001001010101100000",
						 "101010001001010101100110",
						 "101010001001010101101100",
						 "101010001001010101110010",
						 "101010001001010101111000",
						 "101010001001010101111110",
						 "101010001001010110000100",
						 "101010001001010110001010",
						 "101010001001010110010000",
						 "101010001001010110010110",
						 "101010001001010110011100",
						 "101010001001010101000010",
						 "101010001001010101001000",
						 "101010001001010101001110",
						 "101010001001010101010100",
						 "101010001001010101011010",
						 "101010001001010101100000",
						 "101010001001010101100110",
						 "101010001001010101101100",
						 "101010001001010101110010",
						 "101010001001010101111000",
						 "101010001001010101111110",
						 "101010001001010110000100",
						 "101010001001010110001010",
						 "101010001001010110010000",
						 "101010001001010110010110",
						 "101010001001010110011100",
						 "101010001001010101000010",
						 "101010001001010101001000",
						 "101010001001010101001110",
						 "101010001001010101010100",
						 "101010001001010101011010",
						 "101010001001010101100000",
						 "101010001001010101100110",
						 "101010001001010101101100",
						 "101010001001010101110010",
						 "101010001001010101111000",
						 "101010001001010101111110",
						 "101010001001010110000100",
						 "101010001001010110001010",
						 "101010001001010110010000",
						 "101010001001010110010110",
						 "101010001001010110011100",
						 "101010001001010101000010",
						 "101010001001010101000111",
						 "101010001001010101001100",
						 "101010001001010101010001",
						 "101010001001010101010110",
						 "101010001001010101011011",
						 "101010001001010101100000",
						 "101010001001010101100101",
						 "101010001001010101101010",
						 "101010001001010101101111",
						 "101010001001010101110100",
						 "101010001001010101111001",
						 "101010001001010101111110",
						 "101010001001010110000011",
						 "101010001001010110001000",
						 "101010001001010110001101",
						 "101010001001010101000010",
						 "101010001001010101000111",
						 "101010001001010101001100",
						 "101010001001010101010001",
						 "101010001001010101010110",
						 "101010001001010101011011",
						 "101010001001010101100000",
						 "101010001001010101100101",
						 "101010001001010101101010",
						 "101010001001010101101111",
						 "101010001001010101110100",
						 "101010001001010101111001",
						 "101010001001010101111110",
						 "101010001001010110000011",
						 "101010001001010110001000",
						 "101010001001010110001101",
						 "101010001001010101000010",
						 "101010001001010101000110",
						 "101010001001010101001010",
						 "101010001001010101001110",
						 "101010001001010101010010",
						 "101010001001010101010110",
						 "101010001001010101011010",
						 "101010001001010101011110",
						 "101010001001010101100010",
						 "101010001001010101100110",
						 "101010001001010101101010",
						 "101010001001010101101110",
						 "101010001001010101110010",
						 "101010001001010101110110",
						 "101010001001010101111010",
						 "101010001001010101111110",
						 "101010001001010101000010",
						 "101010001001010101000110",
						 "101010001001010101001010",
						 "101010001001010101001110",
						 "101010001001010101010010",
						 "101010001001010101010110",
						 "101010001001010101011010",
						 "101010001001010101011110",
						 "101010001001010101100010",
						 "101010001001010101100110",
						 "101010001001010101101010",
						 "101010001001010101101110",
						 "101010001001010101110010",
						 "101010001001010101110110",
						 "101010001001010101111010",
						 "101010001001010101111110",
						 "101010001001010101000010",
						 "101010001001010101000110",
						 "101010001001010101001010",
						 "101010001001010101001110",
						 "101010001001010101010010",
						 "101010001001010101010110",
						 "101010001001010101011010",
						 "101010001001010101011110",
						 "101010001001010101100010",
						 "101010001001010101100110",
						 "101010001001010101101010",
						 "101010001001010101101110",
						 "101010001001010101110010",
						 "101010001001010101110110",
						 "101010001001010101111010",
						 "101010001001010101111110",
						 "101010001001010101000010",
						 "101010001001010101000101",
						 "101010001001010101001000",
						 "101010001001010101001011",
						 "101010001001010101001110",
						 "101010001001010101010001",
						 "101010001001010101010100",
						 "101010001001010101010111",
						 "101010001001010101011010",
						 "101010001001010101011101",
						 "101010001001010101100000",
						 "101010001001010101100011",
						 "101010001001010101100110",
						 "101010001001010101101001",
						 "101010001001010101101100",
						 "101010001001010101101111",
						 "101010001001010101000010",
						 "101010001001010101000101",
						 "101010001001010101001000",
						 "101010001001010101001011",
						 "101010001001010101001110",
						 "101010001001010101010001",
						 "101010001001010101010100",
						 "101010001001010101010111",
						 "101010001001010101011010",
						 "101010001001010101011101",
						 "101010001001010101100000",
						 "101010001001010101100011",
						 "101010001001010101100110",
						 "101010001001010101101001",
						 "101010001001010101101100",
						 "101010001001010101101111",
						 "101010001001010101000010",
						 "101010001001010101000101",
						 "101010001001010101001000",
						 "101010001001010101001011",
						 "101010001001010101001110",
						 "101010001001010101010001",
						 "101010001001010101010100",
						 "101010001001010101010111",
						 "101010001001010101011010",
						 "101010001001010101011101",
						 "101010001001010101100000",
						 "101010001001010101100011",
						 "101010001001010101100110",
						 "101010001001010101101001",
						 "101010001001010101101100",
						 "101010001001010101101111",
						 "101010001001010101000010",
						 "101010001001010101000100",
						 "101010001001010101000110",
						 "101010001001010101001000",
						 "101010001001010101001010",
						 "101010001001010101001100",
						 "101010001001010101001110",
						 "101010001001010101010000",
						 "101010001001010101010010",
						 "101010001001010101010100",
						 "101010001001010101010110",
						 "101010001001010101011000",
						 "101010001001010101011010",
						 "101010001001010101011100",
						 "101010001001010101011110",
						 "101010001001010101100000",
						 "101010001001010101000010",
						 "101010001001010101000100",
						 "101010001001010101000110",
						 "101010001001010101001000",
						 "101010001001010101001010",
						 "101010001001010101001100",
						 "101010001001010101001110",
						 "101010001001010101010000",
						 "101010001001010101010010",
						 "101010001001010101010100",
						 "101010001001010101010110",
						 "101010001001010101011000",
						 "101010001001010101011010",
						 "101010001001010101011100",
						 "101010001001010101011110",
						 "101010001001010101100000",
						 "101010001001010101000010",
						 "101010001001010101000011",
						 "101010001001010101000100",
						 "101010001001010101000101",
						 "101010001001010101000110",
						 "101010001001010101000111",
						 "101010001001010101001000",
						 "101010001001010101001001",
						 "101010001001010101001010",
						 "101010001001010101001011",
						 "101010001001010101001100",
						 "101010001001010101001101",
						 "101010001001010101001110",
						 "101010001001010101001111",
						 "101010001001010101010000",
						 "101010001001010101010001",
						 "101010001001010101000010",
						 "101010001001010101000011",
						 "101010001001010101000100",
						 "101010001001010101000101",
						 "101010001001010101000110",
						 "101010001001010101000111",
						 "101010001001010101001000",
						 "101010001001010101001001",
						 "101010001001010101001010",
						 "101010001001010101001011",
						 "101010001001010101001100",
						 "101010001001010101001101",
						 "101010001001010101001110",
						 "101010001001010101001111",
						 "101010001001010101010000",
						 "101010001001010101010001",
						 "101010001001010101000010",
						 "101010001001010101000011",
						 "101010001001010101000100",
						 "101010001001010101000101",
						 "101010001001010101000110",
						 "101010001001010101000111",
						 "101010001001010101001000",
						 "101010001001010101001001",
						 "101010001001010101001010",
						 "101010001001010101001011",
						 "101010001001010101001100",
						 "101010001001010101001101",
						 "101010001001010101001110",
						 "101010001001010101001111",
						 "101010001001010101010000",
						 "101010001001010101010001",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101000010",
						 "101010001001010101010001",
						 "101010001001010101010000",
						 "101010001001010101001111",
						 "101010001001010101001110",
						 "101010001001010101001101",
						 "101010001001010101001100",
						 "101010001001010101001011",
						 "101010001001010101001010",
						 "101010001001010101001001",
						 "101010001001010101001000",
						 "101010001001010101000111",
						 "101010001001010101000110",
						 "101010001001010101000101",
						 "101010001001010101000100",
						 "101010001001010101000011",
						 "101010001001010101000010",
						 "101010001001010101010001",
						 "101010001001010101010000",
						 "101010001001010101001111",
						 "101010001001010101001110",
						 "101010001001010101001101",
						 "101010001001010101001100",
						 "101010001001010101001011",
						 "101010001001010101001010",
						 "101010001001010101001001",
						 "101010001001010101001000",
						 "101010001001010101000111",
						 "101010001001010101000110",
						 "101010001001010101000101",
						 "101010001001010101000100",
						 "101010001001010101000011",
						 "101010001001010101000010",
						 "101010001001010101010001",
						 "101010001001010101010000",
						 "101010001001010101001111",
						 "101010001001010101001110",
						 "101010001001010101001101",
						 "101010001001010101001100",
						 "101010001001010101001011",
						 "101010001001010101001010",
						 "101010001001010101001001",
						 "101010001001010101001000",
						 "101010001001010101000111",
						 "101010001001010101000110",
						 "101010001001010101000101",
						 "101010001001010101000100",
						 "101010001001010101000011",
						 "101010001001010101000010",
						 "101010001001010101100000",
						 "101010001001010101011110",
						 "101010001001010101011100",
						 "101010001001010101011010",
						 "101010001001010101011000",
						 "101010001001010101010110",
						 "101010001001010101010100",
						 "101010001001010101010010",
						 "101010001001010101010000",
						 "101010001001010101001110",
						 "101010001001010101001100",
						 "101010001001010101001010",
						 "101010001001010101001000",
						 "101010001001010101000110",
						 "101010001001010101000100",
						 "101010001001010101000010",
						 "101010001001010101100000",
						 "101010001001010101011110",
						 "101010001001010101011100",
						 "101010001001010101011010",
						 "101010001001010101011000",
						 "101010001001010101010110",
						 "101010001001010101010100",
						 "101010001001010101010010",
						 "101010001001010101010000",
						 "101010001001010101001110",
						 "101010001001010101001100",
						 "101010001001010101001010",
						 "101010001001010101001000",
						 "101010001001010101000110",
						 "101010001001010101000100",
						 "101010001001010101000010",
						 "101010001001010101101111",
						 "101010001001010101101100",
						 "101010001001010101101001",
						 "101010001001010101100110",
						 "101010001001010101100011",
						 "101010001001010101100000",
						 "101010001001010101011101",
						 "101010001001010101011010",
						 "101010001001010101010111",
						 "101010001001010101010100",
						 "101010001001010101010001",
						 "101010001001010101001110",
						 "101010001001010101001011",
						 "101010001001010101001000",
						 "101010001001010101000101",
						 "101010001001010101000010",
						 "101010001001010101101111",
						 "101010001001010101101100",
						 "101010001001010101101001",
						 "101010001001010101100110",
						 "101010001001010101100011",
						 "101010001001010101100000",
						 "101010001001010101011101",
						 "101010001001010101011010",
						 "101010001001010101010111",
						 "101010001001010101010100",
						 "101010001001010101010001",
						 "101010001001010101001110",
						 "101010001001010101001011",
						 "101010001001010101001000",
						 "101010001001010101000101",
						 "101010001001010101000010",
						 "101010001001010101101111",
						 "101010001001010101101100",
						 "101010001001010101101001",
						 "101010001001010101100110",
						 "101010001001010101100011",
						 "101010001001010101100000",
						 "101010001001010101011101",
						 "101010001001010101011010",
						 "101010001001010101010111",
						 "101010001001010101010100",
						 "101010001001010101010001",
						 "101010001001010101001110",
						 "101010001001010101001011",
						 "101010001001010101001000",
						 "101010001001010101000101",
						 "101010001001010101000010",
						 "101010001001010101111110",
						 "101010001001010101111010",
						 "101010001001010101110110",
						 "101010001001010101110010",
						 "101010001001010101101110",
						 "101010001001010101101010",
						 "101010001001010101100110",
						 "101010001001010101100010",
						 "101010001001010101011110",
						 "101010001001010101011010",
						 "101010001001010101010110",
						 "101010001001010101010010",
						 "101010001001010101001110",
						 "101010001001010101001010",
						 "101010001001010101000110",
						 "101010001001010101000010",
						 "101010001001010101111110",
						 "101010001001010101111010",
						 "101010001001010101110110",
						 "101010001001010101110010",
						 "101010001001010101101110",
						 "101010001001010101101010",
						 "101010001001010101100110",
						 "101010001001010101100010",
						 "101010001001010101011110",
						 "101010001001010101011010",
						 "101010001001010101010110",
						 "101010001001010101010010",
						 "101010001001010101001110",
						 "101010001001010101001010",
						 "101010001001010101000110",
						 "101010001001010101000010",
						 "101010001001010101111110",
						 "101010001001010101111010",
						 "101010001001010101110110",
						 "101010001001010101110010",
						 "101010001001010101101110",
						 "101010001001010101101010",
						 "101010001001010101100110",
						 "101010001001010101100010",
						 "101010001001010101011110",
						 "101010001001010101011010",
						 "101010001001010101010110",
						 "101010001001010101010010",
						 "101010001001010101001110",
						 "101010001001010101001010",
						 "101010001001010101000110",
						 "101010001001010101000010",
						 "101010001001010110001101",
						 "101010001001010110001000",
						 "101010001001010110000011",
						 "101010001001010101111110",
						 "101010001001010101111001",
						 "101010001001010101110100",
						 "101010001001010101101111",
						 "101010001001010101101010",
						 "101010001001010101100101",
						 "101010001001010101100000",
						 "101010001001010101011011",
						 "101010001001010101010110",
						 "101010001001010101010001",
						 "101010001001010101001100",
						 "101010001001010101000111",
						 "101010001001010101000010",
						 "101010001001010110001101",
						 "101010001001010110001000",
						 "101010001001010110000011",
						 "101010001001010101111110",
						 "101010001001010101111001",
						 "101010001001010101110100",
						 "101010001001010101101111",
						 "101010001001010101101010",
						 "101010001001010101100101",
						 "101010001001010101100000",
						 "101010001001010101011011",
						 "101010001001010101010110",
						 "101010001001010101010001",
						 "101010001001010101001100",
						 "101010001001010101000111",
						 "101010001001010101000010",
						 "101010001001010110011100",
						 "101010001001010110010110",
						 "101010001001010110010000",
						 "101010001001010110001010",
						 "101010001001010110000100",
						 "101010001001010101111110",
						 "101010001001010101111000",
						 "101010001001010101110010",
						 "101010001001010101101100",
						 "101010001001010101100110",
						 "101010001001010101100000",
						 "101010001001010101011010",
						 "101010001001010101010100",
						 "101010001001010101001110",
						 "101010001001010101001000",
						 "101010001001010101000010",
						 "101010001001010110011100",
						 "101010001001010110010110",
						 "101010001001010110010000",
						 "101010001001010110001010",
						 "101010001001010110000100",
						 "101010001001010101111110",
						 "101010001001010101111000",
						 "101010001001010101110010",
						 "101010001001010101101100",
						 "101010001001010101100110",
						 "101010001001010101100000",
						 "101010001001010101011010",
						 "101010001001010101010100",
						 "101010001001010101001110",
						 "101010001001010101001000",
						 "101010001001010101000010",
						 "101010001001010110011100",
						 "101010001001010110010110",
						 "101010001001010110010000",
						 "101010001001010110001010",
						 "101010001001010110000100",
						 "101010001001010101111110",
						 "101010001001010101111000",
						 "101010001001010101110010",
						 "101010001001010101101100",
						 "101010001001010101100110",
						 "101010001001010101100000",
						 "101010001001010101011010",
						 "101010001001010101010100",
						 "101010001001010101001110",
						 "101010001001010101001000",
						 "101010001001010101000010",
						 "101010001001010110101011",
						 "101010001001010110100100",
						 "101010001001010110011101",
						 "101010001001010110010110",
						 "101010001001010110001111",
						 "101010001001010110001000",
						 "101010001001010110000001",
						 "101010001001010101111010",
						 "101010001001010101110011",
						 "101010001001010101101100",
						 "101010001001010101100101",
						 "101010001001010101011110",
						 "101010001001010101010111",
						 "101010001001010101010000",
						 "101010001001010101001001",
						 "101010001001010101000010",
						 "101010001001010110101011",
						 "101010001001010110100100",
						 "101010001001010110011101",
						 "101010001001010110010110",
						 "101010001001010110001111",
						 "101010001001010110001000",
						 "101010001001010110000001",
						 "101010001001010101111010",
						 "101010001001010101110011",
						 "101010001001010101101100",
						 "101010001001010101100101",
						 "101010001001010101011110",
						 "101010001001010101010111",
						 "101010001001010101010000",
						 "101010001001010101001001",
						 "101010001001010101000010",
						 "101010001001010110111010",
						 "101010001001010110110010",
						 "101010001001010110101010",
						 "101010001001010110100010",
						 "101010001001010110011010",
						 "101010001001010110010010",
						 "101010001001010110001010",
						 "101010001001010110000010",
						 "101010001001010101111010",
						 "101010001001010101110010",
						 "101010001001010101101010",
						 "101010001001010101100010",
						 "101010001001010101011010",
						 "101010001001010101010010",
						 "101010001001010101001010",
						 "101010001001010101000010",
						 "101010001001010110111010",
						 "101010001001010110110010",
						 "101010001001010110101010",
						 "101010001001010110100010",
						 "101010001001010110011010",
						 "101010001001010110010010",
						 "101010001001010110001010",
						 "101010001001010110000010",
						 "101010001001010101111010",
						 "101010001001010101110010",
						 "101010001001010101101010",
						 "101010001001010101100010",
						 "101010001001010101011010",
						 "101010001001010101010010",
						 "101010001001010101001010",
						 "101010001001010101000010",
						 "101010001001010110111010",
						 "101010001001010110110010",
						 "101010001001010110101010",
						 "101010001001010110100010",
						 "101010001001010110011010",
						 "101010001001010110010010",
						 "101010001001010110001010",
						 "101010001001010110000010",
						 "101010001001010101111010",
						 "101010001001010101110010",
						 "101010001001010101101010",
						 "101010001001010101100010",
						 "101010001001010101011010",
						 "101010001001010101010010",
						 "101010001001010101001010",
						 "101010001001010101000010",
						 "101010001001010111001001",
						 "101010001001010111000000",
						 "101010001001010110110111",
						 "101010001001010110101110",
						 "101010001001010110100101",
						 "101010001001010110011100",
						 "101010001001010110010011",
						 "101010001001010110001010",
						 "101010001001010110000001",
						 "101010001001010101111000",
						 "101010001001010101101111",
						 "101010001001010101100110",
						 "101010001001010101011101",
						 "101010001001010101010100",
						 "101010001001010101001011",
						 "101010001001010101000010",
						 "101010001001010111001001",
						 "101010001001010111000000",
						 "101010001001010110110111",
						 "101010001001010110101110",
						 "101010001001010110100101",
						 "101010001001010110011100",
						 "101010001001010110010011",
						 "101010001001010110001010",
						 "101010001001010110000001",
						 "101010001001010101111000",
						 "101010001001010101101111",
						 "101010001001010101100110",
						 "101010001001010101011101",
						 "101010001001010101010100",
						 "101010001001010101001011",
						 "101010001001010101000010",
						 "101010001001010111011000",
						 "101010001001010111001110",
						 "101010001001010111000100",
						 "101010001001010110111010",
						 "101010001001010110110000",
						 "101010001001010110100110",
						 "101010001001010110011100",
						 "101010001001010110010010",
						 "101010001001010110001000",
						 "101010001001010101111110",
						 "101010001001010101110100",
						 "101010001001010101101010",
						 "101010001001010101100000",
						 "101010001001010101010110",
						 "101010001001010101001100",
						 "101010001001010101000010",
						 "101010001001010111011000",
						 "101010001001010111001110",
						 "101010001001010111000100",
						 "101010001001010110111010",
						 "101010001001010110110000",
						 "101010001001010110100110",
						 "101010001001010110011100",
						 "101010001001010110010010",
						 "101010001001010110001000",
						 "101010001001010101111110",
						 "101010001001010101110100",
						 "101010001001010101101010",
						 "101010001001010101100000",
						 "101010001001010101010110",
						 "101010001001010101001100",
						 "101010001001010101000010",
						 "101010001001010111011000",
						 "101010001001010111001110",
						 "101010001001010111000100",
						 "101010001001010110111010",
						 "101010001001010110110000",
						 "101010001001010110100110",
						 "101010001001010110011100",
						 "101010001001010110010010",
						 "101010001001010110001000",
						 "101010001001010101111110",
						 "101010001001010101110100",
						 "101010001001010101101010",
						 "101010001001010101100000",
						 "101010001001010101010110",
						 "101010001001010101001100",
						 "101010001001010101000010",
						 "101010001001010111100111",
						 "101010001001010111011100",
						 "101010001001010111010001",
						 "101010001001010111000110",
						 "101010001001010110111011",
						 "101010001001010110110000",
						 "101010001001010110100101",
						 "101010001001010110011010",
						 "101010001001010110001111",
						 "101010001001010110000100",
						 "101010001001010101111001",
						 "101010001001010101101110",
						 "101010001001010101100011",
						 "101010001001010101011000",
						 "101010001001010101001101",
						 "101010001001010101000010",
						 "101010001001010111100111",
						 "101010001001010111011100",
						 "101010001001010111010001",
						 "101010001001010111000110",
						 "101010001001010110111011",
						 "101010001001010110110000",
						 "101010001001010110100101",
						 "101010001001010110011010",
						 "101010001001010110001111",
						 "101010001001010110000100",
						 "101010001001010101111001",
						 "101010001001010101101110",
						 "101010001001010101100011",
						 "101010001001010101011000",
						 "101010001001010101001101",
						 "101010001001010101000010",
						 "101010001001010111110110",
						 "101010001001010111101010",
						 "101010001001010111011110",
						 "101010001001010111010010",
						 "101010001001010111000110",
						 "101010001001010110111010",
						 "101010001001010110101110",
						 "101010001001010110100010",
						 "101010001001010110010110",
						 "101010001001010110001010",
						 "101010001001010101111110",
						 "101010001001010101110010",
						 "101010001001010101100110",
						 "101010001001010101011010",
						 "101010001001010101001110",
						 "101010001001010101000010",
						 "101010001001010111110110",
						 "101010001001010111101010",
						 "101010001001010111011110",
						 "101010001001010111010010",
						 "101010001001010111000110",
						 "101010001001010110111010",
						 "101010001001010110101110",
						 "101010001001010110100010",
						 "101010001001010110010110",
						 "101010001001010110001010",
						 "101010001001010101111110",
						 "101010001001010101110010",
						 "101010001001010101100110",
						 "101010001001010101011010",
						 "101010001001010101001110",
						 "101010001001010101000010",
						 "101010001001010111110110",
						 "101010001001010111101010",
						 "101010001001010111011110",
						 "101010001001010111010010",
						 "101010001001010111000110",
						 "101010001001010110111010",
						 "101010001001010110101110",
						 "101010001001010110100010",
						 "101010001001010110010110",
						 "101010001001010110001010",
						 "101010001001010101111110",
						 "101010001001010101110010",
						 "101010001001010101100110",
						 "101010001001010101011010",
						 "101010001001010101001110",
						 "101010001001010101000010",
						 "101010001001011000000101",
						 "101010001001010111111000",
						 "101010001001010111101011",
						 "101010001001010111011110",
						 "101010001001010111010001",
						 "101010001001010111000100",
						 "101010001001010110110111",
						 "101010001001010110101010",
						 "101010001001010110011101",
						 "101010001001010110010000",
						 "101010001001010110000011",
						 "101010001001010101110110",
						 "101010001001010101101001",
						 "101010001001010101011100",
						 "101010001001010101001111",
						 "101010001001010101000010",
						 "101010001001011000000101",
						 "101010001001010111111000",
						 "101010001001010111101011",
						 "101010001001010111011110",
						 "101010001001010111010001",
						 "101010001001010111000100",
						 "101010001001010110110111",
						 "101010001001010110101010",
						 "101010001001010110011101",
						 "101010001001010110010000",
						 "101010001001010110000011",
						 "101010001001010101110110",
						 "101010001001010101101001",
						 "101010001001010101011100",
						 "101010001001010101001111",
						 "101010001001010101000010",
						 "101010001001011000000101",
						 "101010001001010111111000",
						 "101010001001010111101011",
						 "101010001001010111011110",
						 "101010001001010111010001",
						 "101010001001010111000100",
						 "101010001001010110110111",
						 "101010001001010110101010",
						 "101010001001010110011101",
						 "101010001001010110010000",
						 "101010001001010110000011",
						 "101010001001010101110110",
						 "101010001001010101101001",
						 "101010001001010101011100",
						 "101010001001010101001111",
						 "101010001001010101000010",
						 "101010001001011000010100",
						 "101010001001011000000110",
						 "101010001001010111111000",
						 "101010001001010111101010",
						 "101010001001010111011100",
						 "101010001001010111001110",
						 "101010001001010111000000",
						 "101010001001010110110010",
						 "101010001001010110100100",
						 "101010001001010110010110",
						 "101010001001010110001000",
						 "101010001001010101111010",
						 "101010001001010101101100",
						 "101010001001010101011110",
						 "101010001001010101010000",
						 "101010001001010101000010",
						 "101010001001011000010100",
						 "101010001001011000000110",
						 "101010001001010111111000",
						 "101010001001010111101010",
						 "101010001001010111011100",
						 "101010001001010111001110",
						 "101010001001010111000000",
						 "101010001001010110110010",
						 "101010001001010110100100",
						 "101010001001010110010110",
						 "101010001001010110001000",
						 "101010001001010101111010",
						 "101010001001010101101100",
						 "101010001001010101011110",
						 "101010001001010101010000",
						 "101010001001010101000010",
						 "101010001001011000100011",
						 "101010001001011000010100",
						 "101010001001011000000101",
						 "101010001001010111110110",
						 "101010001001010111100111",
						 "101010001001010111011000",
						 "101010001001010111001001",
						 "101010001001010110111010",
						 "101010001001010110101011",
						 "101010001001010110011100",
						 "101010001001010110001101",
						 "101010001001010101111110",
						 "101010001001010101101111",
						 "101010001001010101100000",
						 "101010001001010101010001",
						 "101010001001010101000010",
						 "101010001001011000100011",
						 "101010001001011000010100",
						 "101010001001011000000101",
						 "101010001001010111110110",
						 "101010001001010111100111",
						 "101010001001010111011000",
						 "101010001001010111001001",
						 "101010001001010110111010",
						 "101010001001010110101011",
						 "101010001001010110011100",
						 "101010001001010110001101",
						 "101010001001010101111110",
						 "101010001001010101101111",
						 "101010001001010101100000",
						 "101010001001010101010001",
						 "101010001001010101000010",
						 "101010001001011000100011",
						 "101010001001011000010100",
						 "101010001001011000000101",
						 "101010001001010111110110",
						 "101010001001010111100111",
						 "101010001001010111011000",
						 "101010001001010111001001",
						 "101010001001010110111010",
						 "101010001001010110101011",
						 "101010001001010110011100",
						 "101010001001010110001101",
						 "101010001001010101111110",
						 "101010001001010101101111",
						 "101010001001010101100000",
						 "101010001001010101010001",
						 "101010001001010101000010",
						 "101010000110110101110100",
						 "101010000110110101100100",
						 "101010000110110101010100",
						 "101010000110110101000100",
						 "101010000110110100110100",
						 "101010000110110100100100",
						 "101010000110110100010100",
						 "101010000110110100000100",
						 "101010000110110011110100",
						 "101010000110110011100100",
						 "101010000110110011010100",
						 "101010000110110011000100",
						 "101010000110110010110100",
						 "101010000110110010100100",
						 "101010000110110010010100",
						 "101010000110110010000100",
						 "101010000110110101110100",
						 "101010000110110101100100",
						 "101010000110110101010100",
						 "101010000110110101000100",
						 "101010000110110100110100",
						 "101010000110110100100100",
						 "101010000110110100010100",
						 "101010000110110100000100",
						 "101010000110110011110100",
						 "101010000110110011100100",
						 "101010000110110011010100",
						 "101010000110110011000100",
						 "101010000110110010110100",
						 "101010000110110010100100",
						 "101010000110110010010100",
						 "101010000110110010000100",
						 "101010000110110110000011",
						 "101010000110110101110010",
						 "101010000110110101100001",
						 "101010000110110101010000",
						 "101010000110110100111111",
						 "101010000110110100101110",
						 "101010000110110100011101",
						 "101010000110110100001100",
						 "101010000110110011111011",
						 "101010000110110011101010",
						 "101010000110110011011001",
						 "101010000110110011001000",
						 "101010000110110010110111",
						 "101010000110110010100110",
						 "101010000110110010010101",
						 "101010000110110010000100",
						 "101010000110110110000011",
						 "101010000110110101110010",
						 "101010000110110101100001",
						 "101010000110110101010000",
						 "101010000110110100111111",
						 "101010000110110100101110",
						 "101010000110110100011101",
						 "101010000110110100001100",
						 "101010000110110011111011",
						 "101010000110110011101010",
						 "101010000110110011011001",
						 "101010000110110011001000",
						 "101010000110110010110111",
						 "101010000110110010100110",
						 "101010000110110010010101",
						 "101010000110110010000100",
						 "101010000110110110000011",
						 "101010000110110101110010",
						 "101010000110110101100001",
						 "101010000110110101010000",
						 "101010000110110100111111",
						 "101010000110110100101110",
						 "101010000110110100011101",
						 "101010000110110100001100",
						 "101010000110110011111011",
						 "101010000110110011101010",
						 "101010000110110011011001",
						 "101010000110110011001000",
						 "101010000110110010110111",
						 "101010000110110010100110",
						 "101010000110110010010101",
						 "101010000110110010000100",
						 "101010000110110110010010",
						 "101010000110110110000000",
						 "101010000110110101101110",
						 "101010000110110101011100",
						 "101010000110110101001010",
						 "101010000110110100111000",
						 "101010000110110100100110",
						 "101010000110110100010100",
						 "101010000110110100000010",
						 "101010000110110011110000",
						 "101010000110110011011110",
						 "101010000110110011001100",
						 "101010000110110010111010",
						 "101010000110110010101000",
						 "101010000110110010010110",
						 "101010000110110010000100",
						 "101010000110110110010010",
						 "101010000110110110000000",
						 "101010000110110101101110",
						 "101010000110110101011100",
						 "101010000110110101001010",
						 "101010000110110100111000",
						 "101010000110110100100110",
						 "101010000110110100010100",
						 "101010000110110100000010",
						 "101010000110110011110000",
						 "101010000110110011011110",
						 "101010000110110011001100",
						 "101010000110110010111010",
						 "101010000110110010101000",
						 "101010000110110010010110",
						 "101010000110110010000100",
						 "101010000110110110100001",
						 "101010000110110110001110",
						 "101010000110110101111011",
						 "101010000110110101101000",
						 "101010000110110101010101",
						 "101010000110110101000010",
						 "101010000110110100101111",
						 "101010000110110100011100",
						 "101010000110110100001001",
						 "101010000110110011110110",
						 "101010000110110011100011",
						 "101010000110110011010000",
						 "101010000110110010111101",
						 "101010000110110010101010",
						 "101010000110110010010111",
						 "101010000110110010000100",
						 "101010000110110110100001",
						 "101010000110110110001110",
						 "101010000110110101111011",
						 "101010000110110101101000",
						 "101010000110110101010101",
						 "101010000110110101000010",
						 "101010000110110100101111",
						 "101010000110110100011100",
						 "101010000110110100001001",
						 "101010000110110011110110",
						 "101010000110110011100011",
						 "101010000110110011010000",
						 "101010000110110010111101",
						 "101010000110110010101010",
						 "101010000110110010010111",
						 "101010000110110010000100",
						 "101010000110110110100001",
						 "101010000110110110001110",
						 "101010000110110101111011",
						 "101010000110110101101000",
						 "101010000110110101010101",
						 "101010000110110101000010",
						 "101010000110110100101111",
						 "101010000110110100011100",
						 "101010000110110100001001",
						 "101010000110110011110110",
						 "101010000110110011100011",
						 "101010000110110011010000",
						 "101010000110110010111101",
						 "101010000110110010101010",
						 "101010000110110010010111",
						 "101010000110110010000100",
						 "101010000110110110110000",
						 "101010000110110110011100",
						 "101010000110110110001000",
						 "101010000110110101110100",
						 "101010000110110101100000",
						 "101010000110110101001100",
						 "101010000110110100111000",
						 "101010000110110100100100",
						 "101010000110110100010000",
						 "101010000110110011111100",
						 "101010000110110011101000",
						 "101010000110110011010100",
						 "101010000110110011000000",
						 "101010000110110010101100",
						 "101010000110110010011000",
						 "101010000110110010000100",
						 "101010000110110110110000",
						 "101010000110110110011100",
						 "101010000110110110001000",
						 "101010000110110101110100",
						 "101010000110110101100000",
						 "101010000110110101001100",
						 "101010000110110100111000",
						 "101010000110110100100100",
						 "101010000110110100010000",
						 "101010000110110011111100",
						 "101010000110110011101000",
						 "101010000110110011010100",
						 "101010000110110011000000",
						 "101010000110110010101100",
						 "101010000110110010011000",
						 "101010000110110010000100",
						 "101010000110110110111111",
						 "101010000110110110101010",
						 "101010000110110110010101",
						 "101010000110110110000000",
						 "101010000110110101101011",
						 "101010000110110101010110",
						 "101010000110110101000001",
						 "101010000110110100101100",
						 "101010000110110100010111",
						 "101010000110110100000010",
						 "101010000110110011101101",
						 "101010000110110011011000",
						 "101010000110110011000011",
						 "101010000110110010101110",
						 "101010000110110010011001",
						 "101010000110110010000100",
						 "101010000110110110111111",
						 "101010000110110110101010",
						 "101010000110110110010101",
						 "101010000110110110000000",
						 "101010000110110101101011",
						 "101010000110110101010110",
						 "101010000110110101000001",
						 "101010000110110100101100",
						 "101010000110110100010111",
						 "101010000110110100000010",
						 "101010000110110011101101",
						 "101010000110110011011000",
						 "101010000110110011000011",
						 "101010000110110010101110",
						 "101010000110110010011001",
						 "101010000110110010000100",
						 "101010000110110110111111",
						 "101010000110110110101010",
						 "101010000110110110010101",
						 "101010000110110110000000",
						 "101010000110110101101011",
						 "101010000110110101010110",
						 "101010000110110101000001",
						 "101010000110110100101100",
						 "101010000110110100010111",
						 "101010000110110100000010",
						 "101010000110110011101101",
						 "101010000110110011011000",
						 "101010000110110011000011",
						 "101010000110110010101110",
						 "101010000110110010011001",
						 "101010000110110010000100",
						 "101010000110110111001110",
						 "101010000110110110111000",
						 "101010000110110110100010",
						 "101010000110110110001100",
						 "101010000110110101110110",
						 "101010000110110101100000",
						 "101010000110110101001010",
						 "101010000110110100110100",
						 "101010000110110100011110",
						 "101010000110110100001000",
						 "101010000110110011110010",
						 "101010000110110011011100",
						 "101010000110110011000110",
						 "101010000110110010110000",
						 "101010000110110010011010",
						 "101010000110110010000100",
						 "101010000110110111001110",
						 "101010000110110110111000",
						 "101010000110110110100010",
						 "101010000110110110001100",
						 "101010000110110101110110",
						 "101010000110110101100000",
						 "101010000110110101001010",
						 "101010000110110100110100",
						 "101010000110110100011110",
						 "101010000110110100001000",
						 "101010000110110011110010",
						 "101010000110110011011100",
						 "101010000110110011000110",
						 "101010000110110010110000",
						 "101010000110110010011010",
						 "101010000110110010000100",
						 "101010000110110111001110",
						 "101010000110110110111000",
						 "101010000110110110100010",
						 "101010000110110110001100",
						 "101010000110110101110110",
						 "101010000110110101100000",
						 "101010000110110101001010",
						 "101010000110110100110100",
						 "101010000110110100011110",
						 "101010000110110100001000",
						 "101010000110110011110010",
						 "101010000110110011011100",
						 "101010000110110011000110",
						 "101010000110110010110000",
						 "101010000110110010011010",
						 "101010000110110010000100",
						 "101010000110110111011101",
						 "101010000110110111000110",
						 "101010000110110110101111",
						 "101010000110110110011000",
						 "101010000110110110000001",
						 "101010000110110101101010",
						 "101010000110110101010011",
						 "101010000110110100111100",
						 "101010000110110100100101",
						 "101010000110110100001110",
						 "101010000110110011110111",
						 "101010000110110011100000",
						 "101010000110110011001001",
						 "101010000110110010110010",
						 "101010000110110010011011",
						 "101010000110110010000100",
						 "101010000110110111011101",
						 "101010000110110111000110",
						 "101010000110110110101111",
						 "101010000110110110011000",
						 "101010000110110110000001",
						 "101010000110110101101010",
						 "101010000110110101010011",
						 "101010000110110100111100",
						 "101010000110110100100101",
						 "101010000110110100001110",
						 "101010000110110011110111",
						 "101010000110110011100000",
						 "101010000110110011001001",
						 "101010000110110010110010",
						 "101010000110110010011011",
						 "101010000110110010000100",
						 "101010000110110111101100",
						 "101010000110110111010100",
						 "101010000110110110111100",
						 "101010000110110110100100",
						 "101010000110110110001100",
						 "101010000110110101110100",
						 "101010000110110101011100",
						 "101010000110110101000100",
						 "101010000110110100101100",
						 "101010000110110100010100",
						 "101010000110110011111100",
						 "101010000110110011100100",
						 "101010000110110011001100",
						 "101010000110110010110100",
						 "101010000110110010011100",
						 "101010000110110010000100",
						 "101010000110110111101100",
						 "101010000110110111010100",
						 "101010000110110110111100",
						 "101010000110110110100100",
						 "101010000110110110001100",
						 "101010000110110101110100",
						 "101010000110110101011100",
						 "101010000110110101000100",
						 "101010000110110100101100",
						 "101010000110110100010100",
						 "101010000110110011111100",
						 "101010000110110011100100",
						 "101010000110110011001100",
						 "101010000110110010110100",
						 "101010000110110010011100",
						 "101010000110110010000100",
						 "101010000110110111101100",
						 "101010000110110111010100",
						 "101010000110110110111100",
						 "101010000110110110100100",
						 "101010000110110110001100",
						 "101010000110110101110100",
						 "101010000110110101011100",
						 "101010000110110101000100",
						 "101010000110110100101100",
						 "101010000110110100010100",
						 "101010000110110011111100",
						 "101010000110110011100100",
						 "101010000110110011001100",
						 "101010000110110010110100",
						 "101010000110110010011100",
						 "101010000110110010000100",
						 "101010000110110111111011",
						 "101010000110110111100010",
						 "101010000110110111001001",
						 "101010000110110110110000",
						 "101010000110110110010111",
						 "101010000110110101111110",
						 "101010000110110101100101",
						 "101010000110110101001100",
						 "101010000110110100110011",
						 "101010000110110100011010",
						 "101010000110110100000001",
						 "101010000110110011101000",
						 "101010000110110011001111",
						 "101010000110110010110110",
						 "101010000110110010011101",
						 "101010000110110010000100",
						 "101010000110110111111011",
						 "101010000110110111100010",
						 "101010000110110111001001",
						 "101010000110110110110000",
						 "101010000110110110010111",
						 "101010000110110101111110",
						 "101010000110110101100101",
						 "101010000110110101001100",
						 "101010000110110100110011",
						 "101010000110110100011010",
						 "101010000110110100000001",
						 "101010000110110011101000",
						 "101010000110110011001111",
						 "101010000110110010110110",
						 "101010000110110010011101",
						 "101010000110110010000100",
						 "101010000110111000001010",
						 "101010000110110111110000",
						 "101010000110110111010110",
						 "101010000110110110111100",
						 "101010000110110110100010",
						 "101010000110110110001000",
						 "101010000110110101101110",
						 "101010000110110101010100",
						 "101010000110110100111010",
						 "101010000110110100100000",
						 "101010000110110100000110",
						 "101010000110110011101100",
						 "101010000110110011010010",
						 "101010000110110010111000",
						 "101010000110110010011110",
						 "101010000110110010000100",
						 "101010000110111000001010",
						 "101010000110110111110000",
						 "101010000110110111010110",
						 "101010000110110110111100",
						 "101010000110110110100010",
						 "101010000110110110001000",
						 "101010000110110101101110",
						 "101010000110110101010100",
						 "101010000110110100111010",
						 "101010000110110100100000",
						 "101010000110110100000110",
						 "101010000110110011101100",
						 "101010000110110011010010",
						 "101010000110110010111000",
						 "101010000110110010011110",
						 "101010000110110010000100",
						 "101010000110111000001010",
						 "101010000110110111110000",
						 "101010000110110111010110",
						 "101010000110110110111100",
						 "101010000110110110100010",
						 "101010000110110110001000",
						 "101010000110110101101110",
						 "101010000110110101010100",
						 "101010000110110100111010",
						 "101010000110110100100000",
						 "101010000110110100000110",
						 "101010000110110011101100",
						 "101010000110110011010010",
						 "101010000110110010111000",
						 "101010000110110010011110",
						 "101010000110110010000100",
						 "101010000110111000011001",
						 "101010000110110111111110",
						 "101010000110110111100011",
						 "101010000110110111001000",
						 "101010000110110110101101",
						 "101010000110110110010010",
						 "101010000110110101110111",
						 "101010000110110101011100",
						 "101010000110110101000001",
						 "101010000110110100100110",
						 "101010000110110100001011",
						 "101010000110110011110000",
						 "101010000110110011010101",
						 "101010000110110010111010",
						 "101010000110110010011111",
						 "101010000110110010000100",
						 "101010000110111000011001",
						 "101010000110110111111110",
						 "101010000110110111100011",
						 "101010000110110111001000",
						 "101010000110110110101101",
						 "101010000110110110010010",
						 "101010000110110101110111",
						 "101010000110110101011100",
						 "101010000110110101000001",
						 "101010000110110100100110",
						 "101010000110110100001011",
						 "101010000110110011110000",
						 "101010000110110011010101",
						 "101010000110110010111010",
						 "101010000110110010011111",
						 "101010000110110010000100",
						 "101010000100010101101010",
						 "101010000100010101001110",
						 "101010000100010100110010",
						 "101010000100010100010110",
						 "101010000100010011111010",
						 "101010000100010011011110",
						 "101010000100010011000010",
						 "101010000100010010100110",
						 "101010000100010010001010",
						 "101010000100010001101110",
						 "101010000100010001010010",
						 "101010000100010000110110",
						 "101010000100010000011010",
						 "101010000100001111111110",
						 "101010000100001111100010",
						 "101010000100001111000110",
						 "101010000100010101101010",
						 "101010000100010101001110",
						 "101010000100010100110010",
						 "101010000100010100010110",
						 "101010000100010011111010",
						 "101010000100010011011110",
						 "101010000100010011000010",
						 "101010000100010010100110",
						 "101010000100010010001010",
						 "101010000100010001101110",
						 "101010000100010001010010",
						 "101010000100010000110110",
						 "101010000100010000011010",
						 "101010000100001111111110",
						 "101010000100001111100010",
						 "101010000100001111000110",
						 "101010000100010101101010",
						 "101010000100010101001110",
						 "101010000100010100110010",
						 "101010000100010100010110",
						 "101010000100010011111010",
						 "101010000100010011011110",
						 "101010000100010011000010",
						 "101010000100010010100110",
						 "101010000100010010001010",
						 "101010000100010001101110",
						 "101010000100010001010010",
						 "101010000100010000110110",
						 "101010000100010000011010",
						 "101010000100001111111110",
						 "101010000100001111100010",
						 "101010000100001111000110",
						 "101010000100010101111001",
						 "101010000100010101011100",
						 "101010000100010100111111",
						 "101010000100010100100010",
						 "101010000100010100000101",
						 "101010000100010011101000",
						 "101010000100010011001011",
						 "101010000100010010101110",
						 "101010000100010010010001",
						 "101010000100010001110100",
						 "101010000100010001010111",
						 "101010000100010000111010",
						 "101010000100010000011101",
						 "101010000100010000000000",
						 "101010000100001111100011",
						 "101010000100001111000110",
						 "101010000100010101111001",
						 "101010000100010101011100",
						 "101010000100010100111111",
						 "101010000100010100100010",
						 "101010000100010100000101",
						 "101010000100010011101000",
						 "101010000100010011001011",
						 "101010000100010010101110",
						 "101010000100010010010001",
						 "101010000100010001110100",
						 "101010000100010001010111",
						 "101010000100010000111010",
						 "101010000100010000011101",
						 "101010000100010000000000",
						 "101010000100001111100011",
						 "101010000100001111000110",
						 "101010000100010101111001",
						 "101010000100010101011100",
						 "101010000100010100111111",
						 "101010000100010100100010",
						 "101010000100010100000101",
						 "101010000100010011101000",
						 "101010000100010011001011",
						 "101010000100010010101110",
						 "101010000100010010010001",
						 "101010000100010001110100",
						 "101010000100010001010111",
						 "101010000100010000111010",
						 "101010000100010000011101",
						 "101010000100010000000000",
						 "101010000100001111100011",
						 "101010000100001111000110",
						 "101010000100010110001000",
						 "101010000100010101101010",
						 "101010000100010101001100",
						 "101010000100010100101110",
						 "101010000100010100010000",
						 "101010000100010011110010",
						 "101010000100010011010100",
						 "101010000100010010110110",
						 "101010000100010010011000",
						 "101010000100010001111010",
						 "101010000100010001011100",
						 "101010000100010000111110",
						 "101010000100010000100000",
						 "101010000100010000000010",
						 "101010000100001111100100",
						 "101010000100001111000110",
						 "101010000100010110001000",
						 "101010000100010101101010",
						 "101010000100010101001100",
						 "101010000100010100101110",
						 "101010000100010100010000",
						 "101010000100010011110010",
						 "101010000100010011010100",
						 "101010000100010010110110",
						 "101010000100010010011000",
						 "101010000100010001111010",
						 "101010000100010001011100",
						 "101010000100010000111110",
						 "101010000100010000100000",
						 "101010000100010000000010",
						 "101010000100001111100100",
						 "101010000100001111000110",
						 "101010000100010110010111",
						 "101010000100010101111000",
						 "101010000100010101011001",
						 "101010000100010100111010",
						 "101010000100010100011011",
						 "101010000100010011111100",
						 "101010000100010011011101",
						 "101010000100010010111110",
						 "101010000100010010011111",
						 "101010000100010010000000",
						 "101010000100010001100001",
						 "101010000100010001000010",
						 "101010000100010000100011",
						 "101010000100010000000100",
						 "101010000100001111100101",
						 "101010000100001111000110",
						 "101010000100010110010111",
						 "101010000100010101111000",
						 "101010000100010101011001",
						 "101010000100010100111010",
						 "101010000100010100011011",
						 "101010000100010011111100",
						 "101010000100010011011101",
						 "101010000100010010111110",
						 "101010000100010010011111",
						 "101010000100010010000000",
						 "101010000100010001100001",
						 "101010000100010001000010",
						 "101010000100010000100011",
						 "101010000100010000000100",
						 "101010000100001111100101",
						 "101010000100001111000110",
						 "101010000100010110010111",
						 "101010000100010101111000",
						 "101010000100010101011001",
						 "101010000100010100111010",
						 "101010000100010100011011",
						 "101010000100010011111100",
						 "101010000100010011011101",
						 "101010000100010010111110",
						 "101010000100010010011111",
						 "101010000100010010000000",
						 "101010000100010001100001",
						 "101010000100010001000010",
						 "101010000100010000100011",
						 "101010000100010000000100",
						 "101010000100001111100101",
						 "101010000100001111000110",
						 "101010000100010110100110",
						 "101010000100010110000110",
						 "101010000100010101100110",
						 "101010000100010101000110",
						 "101010000100010100100110",
						 "101010000100010100000110",
						 "101010000100010011100110",
						 "101010000100010011000110",
						 "101010000100010010100110",
						 "101010000100010010000110",
						 "101010000100010001100110",
						 "101010000100010001000110",
						 "101010000100010000100110",
						 "101010000100010000000110",
						 "101010000100001111100110",
						 "101010000100001111000110",
						 "101010000100010110100110",
						 "101010000100010110000110",
						 "101010000100010101100110",
						 "101010000100010101000110",
						 "101010000100010100100110",
						 "101010000100010100000110",
						 "101010000100010011100110",
						 "101010000100010011000110",
						 "101010000100010010100110",
						 "101010000100010010000110",
						 "101010000100010001100110",
						 "101010000100010001000110",
						 "101010000100010000100110",
						 "101010000100010000000110",
						 "101010000100001111100110",
						 "101010000100001111000110",
						 "101010000100010110110101",
						 "101010000100010110010100",
						 "101010000100010101110011",
						 "101010000100010101010010",
						 "101010000100010100110001",
						 "101010000100010100010000",
						 "101010000100010011101111",
						 "101010000100010011001110",
						 "101010000100010010101101",
						 "101010000100010010001100",
						 "101010000100010001101011",
						 "101010000100010001001010",
						 "101010000100010000101001",
						 "101010000100010000001000",
						 "101010000100001111100111",
						 "101010000100001111000110",
						 "101010000100010110110101",
						 "101010000100010110010100",
						 "101010000100010101110011",
						 "101010000100010101010010",
						 "101010000100010100110001",
						 "101010000100010100010000",
						 "101010000100010011101111",
						 "101010000100010011001110",
						 "101010000100010010101101",
						 "101010000100010010001100",
						 "101010000100010001101011",
						 "101010000100010001001010",
						 "101010000100010000101001",
						 "101010000100010000001000",
						 "101010000100001111100111",
						 "101010000100001111000110",
						 "101010000100010110110101",
						 "101010000100010110010100",
						 "101010000100010101110011",
						 "101010000100010101010010",
						 "101010000100010100110001",
						 "101010000100010100010000",
						 "101010000100010011101111",
						 "101010000100010011001110",
						 "101010000100010010101101",
						 "101010000100010010001100",
						 "101010000100010001101011",
						 "101010000100010001001010",
						 "101010000100010000101001",
						 "101010000100010000001000",
						 "101010000100001111100111",
						 "101010000100001111000110",
						 "101010000100010111000100",
						 "101010000100010110100010",
						 "101010000100010110000000",
						 "101010000100010101011110",
						 "101010000100010100111100",
						 "101010000100010100011010",
						 "101010000100010011111000",
						 "101010000100010011010110",
						 "101010000100010010110100",
						 "101010000100010010010010",
						 "101010000100010001110000",
						 "101010000100010001001110",
						 "101010000100010000101100",
						 "101010000100010000001010",
						 "101010000100001111101000",
						 "101010000100001111000110",
						 "101010000100010111000100",
						 "101010000100010110100010",
						 "101010000100010110000000",
						 "101010000100010101011110",
						 "101010000100010100111100",
						 "101010000100010100011010",
						 "101010000100010011111000",
						 "101010000100010011010110",
						 "101010000100010010110100",
						 "101010000100010010010010",
						 "101010000100010001110000",
						 "101010000100010001001110",
						 "101010000100010000101100",
						 "101010000100010000001010",
						 "101010000100001111101000",
						 "101010000100001111000110",
						 "101010000100010111010011",
						 "101010000100010110110000",
						 "101010000100010110001101",
						 "101010000100010101101010",
						 "101010000100010101000111",
						 "101010000100010100100100",
						 "101010000100010100000001",
						 "101010000100010011011110",
						 "101010000100010010111011",
						 "101010000100010010011000",
						 "101010000100010001110101",
						 "101010000100010001010010",
						 "101010000100010000101111",
						 "101010000100010000001100",
						 "101010000100001111101001",
						 "101010000100001111000110",
						 "101010000100010111010011",
						 "101010000100010110110000",
						 "101010000100010110001101",
						 "101010000100010101101010",
						 "101010000100010101000111",
						 "101010000100010100100100",
						 "101010000100010100000001",
						 "101010000100010011011110",
						 "101010000100010010111011",
						 "101010000100010010011000",
						 "101010000100010001110101",
						 "101010000100010001010010",
						 "101010000100010000101111",
						 "101010000100010000001100",
						 "101010000100001111101001",
						 "101010000100001111000110",
						 "101010000100010111010011",
						 "101010000100010110110000",
						 "101010000100010110001101",
						 "101010000100010101101010",
						 "101010000100010101000111",
						 "101010000100010100100100",
						 "101010000100010100000001",
						 "101010000100010011011110",
						 "101010000100010010111011",
						 "101010000100010010011000",
						 "101010000100010001110101",
						 "101010000100010001010010",
						 "101010000100010000101111",
						 "101010000100010000001100",
						 "101010000100001111101001",
						 "101010000100001111000110",
						 "101010000001110100100100",
						 "101010000001110100000000",
						 "101010000001110011011100",
						 "101010000001110010111000",
						 "101010000001110010010100",
						 "101010000001110001110000",
						 "101010000001110001001100",
						 "101010000001110000101000",
						 "101010000001110000000100",
						 "101010000001101111100000",
						 "101010000001101110111100",
						 "101010000001101110011000",
						 "101010000001101101110100",
						 "101010000001101101010000",
						 "101010000001101100101100",
						 "101010000001101100001000",
						 "101010000001110100100100",
						 "101010000001110100000000",
						 "101010000001110011011100",
						 "101010000001110010111000",
						 "101010000001110010010100",
						 "101010000001110001110000",
						 "101010000001110001001100",
						 "101010000001110000101000",
						 "101010000001110000000100",
						 "101010000001101111100000",
						 "101010000001101110111100",
						 "101010000001101110011000",
						 "101010000001101101110100",
						 "101010000001101101010000",
						 "101010000001101100101100",
						 "101010000001101100001000",
						 "101010000001110100100100",
						 "101010000001110100000000",
						 "101010000001110011011100",
						 "101010000001110010111000",
						 "101010000001110010010100",
						 "101010000001110001110000",
						 "101010000001110001001100",
						 "101010000001110000101000",
						 "101010000001110000000100",
						 "101010000001101111100000",
						 "101010000001101110111100",
						 "101010000001101110011000",
						 "101010000001101101110100",
						 "101010000001101101010000",
						 "101010000001101100101100",
						 "101010000001101100001000",
						 "101010000001110100110011",
						 "101010000001110100001110",
						 "101010000001110011101001",
						 "101010000001110011000100",
						 "101010000001110010011111",
						 "101010000001110001111010",
						 "101010000001110001010101",
						 "101010000001110000110000",
						 "101010000001110000001011",
						 "101010000001101111100110",
						 "101010000001101111000001",
						 "101010000001101110011100",
						 "101010000001101101110111",
						 "101010000001101101010010",
						 "101010000001101100101101",
						 "101010000001101100001000",
						 "101010000001110100110011",
						 "101010000001110100001110",
						 "101010000001110011101001",
						 "101010000001110011000100",
						 "101010000001110010011111",
						 "101010000001110001111010",
						 "101010000001110001010101",
						 "101010000001110000110000",
						 "101010000001110000001011",
						 "101010000001101111100110",
						 "101010000001101111000001",
						 "101010000001101110011100",
						 "101010000001101101110111",
						 "101010000001101101010010",
						 "101010000001101100101101",
						 "101010000001101100001000",
						 "101010000001110101000010",
						 "101010000001110100011100",
						 "101010000001110011110110",
						 "101010000001110011010000",
						 "101010000001110010101010",
						 "101010000001110010000100",
						 "101010000001110001011110",
						 "101010000001110000111000",
						 "101010000001110000010010",
						 "101010000001101111101100",
						 "101010000001101111000110",
						 "101010000001101110100000",
						 "101010000001101101111010",
						 "101010000001101101010100",
						 "101010000001101100101110",
						 "101010000001101100001000",
						 "101010000001110101000010",
						 "101010000001110100011100",
						 "101010000001110011110110",
						 "101010000001110011010000",
						 "101010000001110010101010",
						 "101010000001110010000100",
						 "101010000001110001011110",
						 "101010000001110000111000",
						 "101010000001110000010010",
						 "101010000001101111101100",
						 "101010000001101111000110",
						 "101010000001101110100000",
						 "101010000001101101111010",
						 "101010000001101101010100",
						 "101010000001101100101110",
						 "101010000001101100001000",
						 "101010000001110101000010",
						 "101010000001110100011100",
						 "101010000001110011110110",
						 "101010000001110011010000",
						 "101010000001110010101010",
						 "101010000001110010000100",
						 "101010000001110001011110",
						 "101010000001110000111000",
						 "101010000001110000010010",
						 "101010000001101111101100",
						 "101010000001101111000110",
						 "101010000001101110100000",
						 "101010000001101101111010",
						 "101010000001101101010100",
						 "101010000001101100101110",
						 "101010000001101100001000",
						 "101010000001110101010001",
						 "101010000001110100101010",
						 "101010000001110100000011",
						 "101010000001110011011100",
						 "101010000001110010110101",
						 "101010000001110010001110",
						 "101010000001110001100111",
						 "101010000001110001000000",
						 "101010000001110000011001",
						 "101010000001101111110010",
						 "101010000001101111001011",
						 "101010000001101110100100",
						 "101010000001101101111101",
						 "101010000001101101010110",
						 "101010000001101100101111",
						 "101010000001101100001000",
						 "101010000001110101010001",
						 "101010000001110100101010",
						 "101010000001110100000011",
						 "101010000001110011011100",
						 "101010000001110010110101",
						 "101010000001110010001110",
						 "101010000001110001100111",
						 "101010000001110001000000",
						 "101010000001110000011001",
						 "101010000001101111110010",
						 "101010000001101111001011",
						 "101010000001101110100100",
						 "101010000001101101111101",
						 "101010000001101101010110",
						 "101010000001101100101111",
						 "101010000001101100001000",
						 "101010000001110101100000",
						 "101010000001110100111000",
						 "101010000001110100010000",
						 "101010000001110011101000",
						 "101010000001110011000000",
						 "101010000001110010011000",
						 "101010000001110001110000",
						 "101010000001110001001000",
						 "101010000001110000100000",
						 "101010000001101111111000",
						 "101010000001101111010000",
						 "101010000001101110101000",
						 "101010000001101110000000",
						 "101010000001101101011000",
						 "101010000001101100110000",
						 "101010000001101100001000",
						 "101010000001110101100000",
						 "101010000001110100111000",
						 "101010000001110100010000",
						 "101010000001110011101000",
						 "101010000001110011000000",
						 "101010000001110010011000",
						 "101010000001110001110000",
						 "101010000001110001001000",
						 "101010000001110000100000",
						 "101010000001101111111000",
						 "101010000001101111010000",
						 "101010000001101110101000",
						 "101010000001101110000000",
						 "101010000001101101011000",
						 "101010000001101100110000",
						 "101010000001101100001000",
						 "101010000001110101100000",
						 "101010000001110100111000",
						 "101010000001110100010000",
						 "101010000001110011101000",
						 "101010000001110011000000",
						 "101010000001110010011000",
						 "101010000001110001110000",
						 "101010000001110001001000",
						 "101010000001110000100000",
						 "101010000001101111111000",
						 "101010000001101111010000",
						 "101010000001101110101000",
						 "101010000001101110000000",
						 "101010000001101101011000",
						 "101010000001101100110000",
						 "101010000001101100001000",
						 "101010000001110101101111",
						 "101010000001110101000110",
						 "101010000001110100011101",
						 "101010000001110011110100",
						 "101010000001110011001011",
						 "101010000001110010100010",
						 "101010000001110001111001",
						 "101010000001110001010000",
						 "101010000001110000100111",
						 "101010000001101111111110",
						 "101010000001101111010101",
						 "101010000001101110101100",
						 "101010000001101110000011",
						 "101010000001101101011010",
						 "101010000001101100110001",
						 "101010000001101100001000",
						 "101010000001110101101111",
						 "101010000001110101000110",
						 "101010000001110100011101",
						 "101010000001110011110100",
						 "101010000001110011001011",
						 "101010000001110010100010",
						 "101010000001110001111001",
						 "101010000001110001010000",
						 "101010000001110000100111",
						 "101010000001101111111110",
						 "101010000001101111010101",
						 "101010000001101110101100",
						 "101010000001101110000011",
						 "101010000001101101011010",
						 "101010000001101100110001",
						 "101010000001101100001000",
						 "101010000001110101101111",
						 "101010000001110101000110",
						 "101010000001110100011101",
						 "101010000001110011110100",
						 "101010000001110011001011",
						 "101010000001110010100010",
						 "101010000001110001111001",
						 "101010000001110001010000",
						 "101010000001110000100111",
						 "101010000001101111111110",
						 "101010000001101111010101",
						 "101010000001101110101100",
						 "101010000001101110000011",
						 "101010000001101101011010",
						 "101010000001101100110001",
						 "101010000001101100001000",
						 "101010000001110101111110",
						 "101010000001110101010100",
						 "101010000001110100101010",
						 "101010000001110100000000",
						 "101010000001110011010110",
						 "101010000001110010101100",
						 "101010000001110010000010",
						 "101010000001110001011000",
						 "101010000001110000101110",
						 "101010000001110000000100",
						 "101010000001101111011010",
						 "101010000001101110110000",
						 "101010000001101110000110",
						 "101010000001101101011100",
						 "101010000001101100110010",
						 "101010000001101100001000",
						 "101001111111010011000000",
						 "101001111111010010010110",
						 "101001111111010001101100",
						 "101001111111010001000010",
						 "101001111111010000011000",
						 "101001111111001111101110",
						 "101001111111001111000100",
						 "101001111111001110011010",
						 "101001111111001101110000",
						 "101001111111001101000110",
						 "101001111111001100011100",
						 "101001111111001011110010",
						 "101001111111001011001000",
						 "101001111111001010011110",
						 "101001111111001001110100",
						 "101001111111001001001010",
						 "101001111111010011001111",
						 "101001111111010010100100",
						 "101001111111010001111001",
						 "101001111111010001001110",
						 "101001111111010000100011",
						 "101001111111001111111000",
						 "101001111111001111001101",
						 "101001111111001110100010",
						 "101001111111001101110111",
						 "101001111111001101001100",
						 "101001111111001100100001",
						 "101001111111001011110110",
						 "101001111111001011001011",
						 "101001111111001010100000",
						 "101001111111001001110101",
						 "101001111111001001001010",
						 "101001111111010011001111",
						 "101001111111010010100100",
						 "101001111111010001111001",
						 "101001111111010001001110",
						 "101001111111010000100011",
						 "101001111111001111111000",
						 "101001111111001111001101",
						 "101001111111001110100010",
						 "101001111111001101110111",
						 "101001111111001101001100",
						 "101001111111001100100001",
						 "101001111111001011110110",
						 "101001111111001011001011",
						 "101001111111001010100000",
						 "101001111111001001110101",
						 "101001111111001001001010",
						 "101001111111010011001111",
						 "101001111111010010100100",
						 "101001111111010001111001",
						 "101001111111010001001110",
						 "101001111111010000100011",
						 "101001111111001111111000",
						 "101001111111001111001101",
						 "101001111111001110100010",
						 "101001111111001101110111",
						 "101001111111001101001100",
						 "101001111111001100100001",
						 "101001111111001011110110",
						 "101001111111001011001011",
						 "101001111111001010100000",
						 "101001111111001001110101",
						 "101001111111001001001010",
						 "101001111111010011011110",
						 "101001111111010010110010",
						 "101001111111010010000110",
						 "101001111111010001011010",
						 "101001111111010000101110",
						 "101001111111010000000010",
						 "101001111111001111010110",
						 "101001111111001110101010",
						 "101001111111001101111110",
						 "101001111111001101010010",
						 "101001111111001100100110",
						 "101001111111001011111010",
						 "101001111111001011001110",
						 "101001111111001010100010",
						 "101001111111001001110110",
						 "101001111111001001001010",
						 "101001111111010011011110",
						 "101001111111010010110010",
						 "101001111111010010000110",
						 "101001111111010001011010",
						 "101001111111010000101110",
						 "101001111111010000000010",
						 "101001111111001111010110",
						 "101001111111001110101010",
						 "101001111111001101111110",
						 "101001111111001101010010",
						 "101001111111001100100110",
						 "101001111111001011111010",
						 "101001111111001011001110",
						 "101001111111001010100010",
						 "101001111111001001110110",
						 "101001111111001001001010",
						 "101001111111010011101101",
						 "101001111111010011000000",
						 "101001111111010010010011",
						 "101001111111010001100110",
						 "101001111111010000111001",
						 "101001111111010000001100",
						 "101001111111001111011111",
						 "101001111111001110110010",
						 "101001111111001110000101",
						 "101001111111001101011000",
						 "101001111111001100101011",
						 "101001111111001011111110",
						 "101001111111001011010001",
						 "101001111111001010100100",
						 "101001111111001001110111",
						 "101001111111001001001010",
						 "101001111111010011101101",
						 "101001111111010011000000",
						 "101001111111010010010011",
						 "101001111111010001100110",
						 "101001111111010000111001",
						 "101001111111010000001100",
						 "101001111111001111011111",
						 "101001111111001110110010",
						 "101001111111001110000101",
						 "101001111111001101011000",
						 "101001111111001100101011",
						 "101001111111001011111110",
						 "101001111111001011010001",
						 "101001111111001010100100",
						 "101001111111001001110111",
						 "101001111111001001001010",
						 "101001111111010011101101",
						 "101001111111010011000000",
						 "101001111111010010010011",
						 "101001111111010001100110",
						 "101001111111010000111001",
						 "101001111111010000001100",
						 "101001111111001111011111",
						 "101001111111001110110010",
						 "101001111111001110000101",
						 "101001111111001101011000",
						 "101001111111001100101011",
						 "101001111111001011111110",
						 "101001111111001011010001",
						 "101001111111001010100100",
						 "101001111111001001110111",
						 "101001111111001001001010",
						 "101001111111010011111100",
						 "101001111111010011001110",
						 "101001111111010010100000",
						 "101001111111010001110010",
						 "101001111111010001000100",
						 "101001111111010000010110",
						 "101001111111001111101000",
						 "101001111111001110111010",
						 "101001111111001110001100",
						 "101001111111001101011110",
						 "101001111111001100110000",
						 "101001111111001100000010",
						 "101001111111001011010100",
						 "101001111111001010100110",
						 "101001111111001001111000",
						 "101001111111001001001010",
						 "101001111111010011111100",
						 "101001111111010011001110",
						 "101001111111010010100000",
						 "101001111111010001110010",
						 "101001111111010001000100",
						 "101001111111010000010110",
						 "101001111111001111101000",
						 "101001111111001110111010",
						 "101001111111001110001100",
						 "101001111111001101011110",
						 "101001111111001100110000",
						 "101001111111001100000010",
						 "101001111111001011010100",
						 "101001111111001010100110",
						 "101001111111001001111000",
						 "101001111111001001001010",
						 "101001111111010011111100",
						 "101001111111010011001110",
						 "101001111111010010100000",
						 "101001111111010001110010",
						 "101001111111010001000100",
						 "101001111111010000010110",
						 "101001111111001111101000",
						 "101001111111001110111010",
						 "101001111111001110001100",
						 "101001111111001101011110",
						 "101001111111001100110000",
						 "101001111111001100000010",
						 "101001111111001011010100",
						 "101001111111001010100110",
						 "101001111111001001111000",
						 "101001111111001001001010",
						 "101001111111010100001011",
						 "101001111111010011011100",
						 "101001111111010010101101",
						 "101001111111010001111110",
						 "101001111111010001001111",
						 "101001111111010000100000",
						 "101001111111001111110001",
						 "101001111111001111000010",
						 "101001111111001110010011",
						 "101001111111001101100100",
						 "101001111111001100110101",
						 "101001111111001100000110",
						 "101001111111001011010111",
						 "101001111111001010101000",
						 "101001111111001001111001",
						 "101001111111001001001010",
						 "101001111111010100001011",
						 "101001111111010011011100",
						 "101001111111010010101101",
						 "101001111111010001111110",
						 "101001111111010001001111",
						 "101001111111010000100000",
						 "101001111111001111110001",
						 "101001111111001111000010",
						 "101001111111001110010011",
						 "101001111111001101100100",
						 "101001111111001100110101",
						 "101001111111001100000110",
						 "101001111111001011010111",
						 "101001111111001010101000",
						 "101001111111001001111001",
						 "101001111111001001001010",
						 "101001111100110001011100",
						 "101001111100110000101100",
						 "101001111100101111111100",
						 "101001111100101111001100",
						 "101001111100101110011100",
						 "101001111100101101101100",
						 "101001111100101100111100",
						 "101001111100101100001100",
						 "101001111100101011011100",
						 "101001111100101010101100",
						 "101001111100101001111100",
						 "101001111100101001001100",
						 "101001111100101000011100",
						 "101001111100100111101100",
						 "101001111100100110111100",
						 "101001111100100110001100",
						 "101001111100110001011100",
						 "101001111100110000101100",
						 "101001111100101111111100",
						 "101001111100101111001100",
						 "101001111100101110011100",
						 "101001111100101101101100",
						 "101001111100101100111100",
						 "101001111100101100001100",
						 "101001111100101011011100",
						 "101001111100101010101100",
						 "101001111100101001111100",
						 "101001111100101001001100",
						 "101001111100101000011100",
						 "101001111100100111101100",
						 "101001111100100110111100",
						 "101001111100100110001100",
						 "101001111100110001011100",
						 "101001111100110000101100",
						 "101001111100101111111100",
						 "101001111100101111001100",
						 "101001111100101110011100",
						 "101001111100101101101100",
						 "101001111100101100111100",
						 "101001111100101100001100",
						 "101001111100101011011100",
						 "101001111100101010101100",
						 "101001111100101001111100",
						 "101001111100101001001100",
						 "101001111100101000011100",
						 "101001111100100111101100",
						 "101001111100100110111100",
						 "101001111100100110001100",
						 "101001111100110001101011",
						 "101001111100110000111010",
						 "101001111100110000001001",
						 "101001111100101111011000",
						 "101001111100101110100111",
						 "101001111100101101110110",
						 "101001111100101101000101",
						 "101001111100101100010100",
						 "101001111100101011100011",
						 "101001111100101010110010",
						 "101001111100101010000001",
						 "101001111100101001010000",
						 "101001111100101000011111",
						 "101001111100100111101110",
						 "101001111100100110111101",
						 "101001111100100110001100",
						 "101001111100110001101011",
						 "101001111100110000111010",
						 "101001111100110000001001",
						 "101001111100101111011000",
						 "101001111100101110100111",
						 "101001111100101101110110",
						 "101001111100101101000101",
						 "101001111100101100010100",
						 "101001111100101011100011",
						 "101001111100101010110010",
						 "101001111100101010000001",
						 "101001111100101001010000",
						 "101001111100101000011111",
						 "101001111100100111101110",
						 "101001111100100110111101",
						 "101001111100100110001100",
						 "101001111100110001111010",
						 "101001111100110001001000",
						 "101001111100110000010110",
						 "101001111100101111100100",
						 "101001111100101110110010",
						 "101001111100101110000000",
						 "101001111100101101001110",
						 "101001111100101100011100",
						 "101001111100101011101010",
						 "101001111100101010111000",
						 "101001111100101010000110",
						 "101001111100101001010100",
						 "101001111100101000100010",
						 "101001111100100111110000",
						 "101001111100100110111110",
						 "101001111100100110001100",
						 "101001111100110001111010",
						 "101001111100110001001000",
						 "101001111100110000010110",
						 "101001111100101111100100",
						 "101001111100101110110010",
						 "101001111100101110000000",
						 "101001111100101101001110",
						 "101001111100101100011100",
						 "101001111100101011101010",
						 "101001111100101010111000",
						 "101001111100101010000110",
						 "101001111100101001010100",
						 "101001111100101000100010",
						 "101001111100100111110000",
						 "101001111100100110111110",
						 "101001111100100110001100",
						 "101001111100110001111010",
						 "101001111100110001001000",
						 "101001111100110000010110",
						 "101001111100101111100100",
						 "101001111100101110110010",
						 "101001111100101110000000",
						 "101001111100101101001110",
						 "101001111100101100011100",
						 "101001111100101011101010",
						 "101001111100101010111000",
						 "101001111100101010000110",
						 "101001111100101001010100",
						 "101001111100101000100010",
						 "101001111100100111110000",
						 "101001111100100110111110",
						 "101001111100100110001100",
						 "101001111100110010001001",
						 "101001111100110001010110",
						 "101001111100110000100011",
						 "101001111100101111110000",
						 "101001111100101110111101",
						 "101001111100101110001010",
						 "101001111100101101010111",
						 "101001111100101100100100",
						 "101001111100101011110001",
						 "101001111100101010111110",
						 "101001111100101010001011",
						 "101001111100101001011000",
						 "101001111100101000100101",
						 "101001111100100111110010",
						 "101001111100100110111111",
						 "101001111100100110001100",
						 "101001111100110010001001",
						 "101001111100110001010110",
						 "101001111100110000100011",
						 "101001111100101111110000",
						 "101001111100101110111101",
						 "101001111100101110001010",
						 "101001111100101101010111",
						 "101001111100101100100100",
						 "101001111100101011110001",
						 "101001111100101010111110",
						 "101001111100101010001011",
						 "101001111100101001011000",
						 "101001111100101000100101",
						 "101001111100100111110010",
						 "101001111100100110111111",
						 "101001111100100110001100",
						 "101001111100110010001001",
						 "101001111100110001010110",
						 "101001111100110000100011",
						 "101001111100101111110000",
						 "101001111100101110111101",
						 "101001111100101110001010",
						 "101001111100101101010111",
						 "101001111100101100100100",
						 "101001111100101011110001",
						 "101001111100101010111110",
						 "101001111100101010001011",
						 "101001111100101001011000",
						 "101001111100101000100101",
						 "101001111100100111110010",
						 "101001111100100110111111",
						 "101001111100100110001100",
						 "101001111100110010011000",
						 "101001111100110001100100",
						 "101001111100110000110000",
						 "101001111100101111111100",
						 "101001111100101111001000",
						 "101001111100101110010100",
						 "101001111100101101100000",
						 "101001111100101100101100",
						 "101001111100101011111000",
						 "101001111100101011000100",
						 "101001111100101010010000",
						 "101001111100101001011100",
						 "101001111100101000101000",
						 "101001111100100111110100",
						 "101001111100100111000000",
						 "101001111100100110001100",
						 "101001111100110010011000",
						 "101001111100110001100100",
						 "101001111100110000110000",
						 "101001111100101111111100",
						 "101001111100101111001000",
						 "101001111100101110010100",
						 "101001111100101101100000",
						 "101001111100101100101100",
						 "101001111100101011111000",
						 "101001111100101011000100",
						 "101001111100101010010000",
						 "101001111100101001011100",
						 "101001111100101000101000",
						 "101001111100100111110100",
						 "101001111100100111000000",
						 "101001111100100110001100",
						 "101001111010001111101001",
						 "101001111010001110110100",
						 "101001111010001101111111",
						 "101001111010001101001010",
						 "101001111010001100010101",
						 "101001111010001011100000",
						 "101001111010001010101011",
						 "101001111010001001110110",
						 "101001111010001001000001",
						 "101001111010001000001100",
						 "101001111010000111010111",
						 "101001111010000110100010",
						 "101001111010000101101101",
						 "101001111010000100111000",
						 "101001111010000100000011",
						 "101001111010000011001110",
						 "101001111010001111101001",
						 "101001111010001110110100",
						 "101001111010001101111111",
						 "101001111010001101001010",
						 "101001111010001100010101",
						 "101001111010001011100000",
						 "101001111010001010101011",
						 "101001111010001001110110",
						 "101001111010001001000001",
						 "101001111010001000001100",
						 "101001111010000111010111",
						 "101001111010000110100010",
						 "101001111010000101101101",
						 "101001111010000100111000",
						 "101001111010000100000011",
						 "101001111010000011001110",
						 "101001111010001111101001",
						 "101001111010001110110100",
						 "101001111010001101111111",
						 "101001111010001101001010",
						 "101001111010001100010101",
						 "101001111010001011100000",
						 "101001111010001010101011",
						 "101001111010001001110110",
						 "101001111010001001000001",
						 "101001111010001000001100",
						 "101001111010000111010111",
						 "101001111010000110100010",
						 "101001111010000101101101",
						 "101001111010000100111000",
						 "101001111010000100000011",
						 "101001111010000011001110",
						 "101001111010001111111000",
						 "101001111010001111000010",
						 "101001111010001110001100",
						 "101001111010001101010110",
						 "101001111010001100100000",
						 "101001111010001011101010",
						 "101001111010001010110100",
						 "101001111010001001111110",
						 "101001111010001001001000",
						 "101001111010001000010010",
						 "101001111010000111011100",
						 "101001111010000110100110",
						 "101001111010000101110000",
						 "101001111010000100111010",
						 "101001111010000100000100",
						 "101001111010000011001110",
						 "101001111010001111111000",
						 "101001111010001111000010",
						 "101001111010001110001100",
						 "101001111010001101010110",
						 "101001111010001100100000",
						 "101001111010001011101010",
						 "101001111010001010110100",
						 "101001111010001001111110",
						 "101001111010001001001000",
						 "101001111010001000010010",
						 "101001111010000111011100",
						 "101001111010000110100110",
						 "101001111010000101110000",
						 "101001111010000100111010",
						 "101001111010000100000100",
						 "101001111010000011001110",
						 "101001111010010000000111",
						 "101001111010001111010000",
						 "101001111010001110011001",
						 "101001111010001101100010",
						 "101001111010001100101011",
						 "101001111010001011110100",
						 "101001111010001010111101",
						 "101001111010001010000110",
						 "101001111010001001001111",
						 "101001111010001000011000",
						 "101001111010000111100001",
						 "101001111010000110101010",
						 "101001111010000101110011",
						 "101001111010000100111100",
						 "101001111010000100000101",
						 "101001111010000011001110",
						 "101001111010010000000111",
						 "101001111010001111010000",
						 "101001111010001110011001",
						 "101001111010001101100010",
						 "101001111010001100101011",
						 "101001111010001011110100",
						 "101001111010001010111101",
						 "101001111010001010000110",
						 "101001111010001001001111",
						 "101001111010001000011000",
						 "101001111010000111100001",
						 "101001111010000110101010",
						 "101001111010000101110011",
						 "101001111010000100111100",
						 "101001111010000100000101",
						 "101001111010000011001110",
						 "101001111010010000000111",
						 "101001111010001111010000",
						 "101001111010001110011001",
						 "101001111010001101100010",
						 "101001111010001100101011",
						 "101001111010001011110100",
						 "101001111010001010111101",
						 "101001111010001010000110",
						 "101001111010001001001111",
						 "101001111010001000011000",
						 "101001111010000111100001",
						 "101001111010000110101010",
						 "101001111010000101110011",
						 "101001111010000100111100",
						 "101001111010000100000101",
						 "101001111010000011001110",
						 "101001111010010000010110",
						 "101001111010001111011110",
						 "101001111010001110100110",
						 "101001111010001101101110",
						 "101001111010001100110110",
						 "101001111010001011111110",
						 "101001111010001011000110",
						 "101001111010001010001110",
						 "101001111010001001010110",
						 "101001111010001000011110",
						 "101001111010000111100110",
						 "101001111010000110101110",
						 "101001111010000101110110",
						 "101001111010000100111110",
						 "101001111010000100000110",
						 "101001111010000011001110",
						 "101001111010010000010110",
						 "101001111010001111011110",
						 "101001111010001110100110",
						 "101001111010001101101110",
						 "101001111010001100110110",
						 "101001111010001011111110",
						 "101001111010001011000110",
						 "101001111010001010001110",
						 "101001111010001001010110",
						 "101001111010001000011110",
						 "101001111010000111100110",
						 "101001111010000110101110",
						 "101001111010000101110110",
						 "101001111010000100111110",
						 "101001111010000100000110",
						 "101001111010000011001110",
						 "101001111010010000010110",
						 "101001111010001111011110",
						 "101001111010001110100110",
						 "101001111010001101101110",
						 "101001111010001100110110",
						 "101001111010001011111110",
						 "101001111010001011000110",
						 "101001111010001010001110",
						 "101001111010001001010110",
						 "101001111010001000011110",
						 "101001111010000111100110",
						 "101001111010000110101110",
						 "101001111010000101110110",
						 "101001111010000100111110",
						 "101001111010000100000110",
						 "101001111010000011001110",
						 "101001111010010000100101",
						 "101001111010001111101100",
						 "101001111010001110110011",
						 "101001111010001101111010",
						 "101001111010001101000001",
						 "101001111010001100001000",
						 "101001111010001011001111",
						 "101001111010001010010110",
						 "101001111010001001011101",
						 "101001111010001000100100",
						 "101001111010000111101011",
						 "101001111010000110110010",
						 "101001111010000101111001",
						 "101001111010000101000000",
						 "101001111010000100000111",
						 "101001111010000011001110",
						 "101001110111101101100111",
						 "101001110111101100101110",
						 "101001110111101011110101",
						 "101001110111101010111100",
						 "101001110111101010000011",
						 "101001110111101001001010",
						 "101001110111101000010001",
						 "101001110111100111011000",
						 "101001110111100110011111",
						 "101001110111100101100110",
						 "101001110111100100101101",
						 "101001110111100011110100",
						 "101001110111100010111011",
						 "101001110111100010000010",
						 "101001110111100001001001",
						 "101001110111100000010000",
						 "101001110111101101110110",
						 "101001110111101100111100",
						 "101001110111101100000010",
						 "101001110111101011001000",
						 "101001110111101010001110",
						 "101001110111101001010100",
						 "101001110111101000011010",
						 "101001110111100111100000",
						 "101001110111100110100110",
						 "101001110111100101101100",
						 "101001110111100100110010",
						 "101001110111100011111000",
						 "101001110111100010111110",
						 "101001110111100010000100",
						 "101001110111100001001010",
						 "101001110111100000010000",
						 "101001110111101101110110",
						 "101001110111101100111100",
						 "101001110111101100000010",
						 "101001110111101011001000",
						 "101001110111101010001110",
						 "101001110111101001010100",
						 "101001110111101000011010",
						 "101001110111100111100000",
						 "101001110111100110100110",
						 "101001110111100101101100",
						 "101001110111100100110010",
						 "101001110111100011111000",
						 "101001110111100010111110",
						 "101001110111100010000100",
						 "101001110111100001001010",
						 "101001110111100000010000",
						 "101001110111101101110110",
						 "101001110111101100111100",
						 "101001110111101100000010",
						 "101001110111101011001000",
						 "101001110111101010001110",
						 "101001110111101001010100",
						 "101001110111101000011010",
						 "101001110111100111100000",
						 "101001110111100110100110",
						 "101001110111100101101100",
						 "101001110111100100110010",
						 "101001110111100011111000",
						 "101001110111100010111110",
						 "101001110111100010000100",
						 "101001110111100001001010",
						 "101001110111100000010000",
						 "101001110111101110000101",
						 "101001110111101101001010",
						 "101001110111101100001111",
						 "101001110111101011010100",
						 "101001110111101010011001",
						 "101001110111101001011110",
						 "101001110111101000100011",
						 "101001110111100111101000",
						 "101001110111100110101101",
						 "101001110111100101110010",
						 "101001110111100100110111",
						 "101001110111100011111100",
						 "101001110111100011000001",
						 "101001110111100010000110",
						 "101001110111100001001011",
						 "101001110111100000010000",
						 "101001110111101110000101",
						 "101001110111101101001010",
						 "101001110111101100001111",
						 "101001110111101011010100",
						 "101001110111101010011001",
						 "101001110111101001011110",
						 "101001110111101000100011",
						 "101001110111100111101000",
						 "101001110111100110101101",
						 "101001110111100101110010",
						 "101001110111100100110111",
						 "101001110111100011111100",
						 "101001110111100011000001",
						 "101001110111100010000110",
						 "101001110111100001001011",
						 "101001110111100000010000",
						 "101001110111101110000101",
						 "101001110111101101001010",
						 "101001110111101100001111",
						 "101001110111101011010100",
						 "101001110111101010011001",
						 "101001110111101001011110",
						 "101001110111101000100011",
						 "101001110111100111101000",
						 "101001110111100110101101",
						 "101001110111100101110010",
						 "101001110111100100110111",
						 "101001110111100011111100",
						 "101001110111100011000001",
						 "101001110111100010000110",
						 "101001110111100001001011",
						 "101001110111100000010000",
						 "101001110111101110010100",
						 "101001110111101101011000",
						 "101001110111101100011100",
						 "101001110111101011100000",
						 "101001110111101010100100",
						 "101001110111101001101000",
						 "101001110111101000101100",
						 "101001110111100111110000",
						 "101001110111100110110100",
						 "101001110111100101111000",
						 "101001110111100100111100",
						 "101001110111100100000000",
						 "101001110111100011000100",
						 "101001110111100010001000",
						 "101001110111100001001100",
						 "101001110111100000010000",
						 "101001110111101110010100",
						 "101001110111101101011000",
						 "101001110111101100011100",
						 "101001110111101011100000",
						 "101001110111101010100100",
						 "101001110111101001101000",
						 "101001110111101000101100",
						 "101001110111100111110000",
						 "101001110111100110110100",
						 "101001110111100101111000",
						 "101001110111100100111100",
						 "101001110111100100000000",
						 "101001110111100011000100",
						 "101001110111100010001000",
						 "101001110111100001001100",
						 "101001110111100000010000",
						 "101001110111101110100011",
						 "101001110111101101100110",
						 "101001110111101100101001",
						 "101001110111101011101100",
						 "101001110111101010101111",
						 "101001110111101001110010",
						 "101001110111101000110101",
						 "101001110111100111111000",
						 "101001110111100110111011",
						 "101001110111100101111110",
						 "101001110111100101000001",
						 "101001110111100100000100",
						 "101001110111100011000111",
						 "101001110111100010001010",
						 "101001110111100001001101",
						 "101001110111100000010000",
						 "101001110111101110100011",
						 "101001110111101101100110",
						 "101001110111101100101001",
						 "101001110111101011101100",
						 "101001110111101010101111",
						 "101001110111101001110010",
						 "101001110111101000110101",
						 "101001110111100111111000",
						 "101001110111100110111011",
						 "101001110111100101111110",
						 "101001110111100101000001",
						 "101001110111100100000100",
						 "101001110111100011000111",
						 "101001110111100010001010",
						 "101001110111100001001101",
						 "101001110111100000010000",
						 "101001110101001011100101",
						 "101001110101001010101000",
						 "101001110101001001101011",
						 "101001110101001000101110",
						 "101001110101000111110001",
						 "101001110101000110110100",
						 "101001110101000101110111",
						 "101001110101000100111010",
						 "101001110101000011111101",
						 "101001110101000011000000",
						 "101001110101000010000011",
						 "101001110101000001000110",
						 "101001110101000000001001",
						 "101001110100111111001100",
						 "101001110100111110001111",
						 "101001110100111101010010",
						 "101001110101001011110100",
						 "101001110101001010110110",
						 "101001110101001001111000",
						 "101001110101001000111010",
						 "101001110101000111111100",
						 "101001110101000110111110",
						 "101001110101000110000000",
						 "101001110101000101000010",
						 "101001110101000100000100",
						 "101001110101000011000110",
						 "101001110101000010001000",
						 "101001110101000001001010",
						 "101001110101000000001100",
						 "101001110100111111001110",
						 "101001110100111110010000",
						 "101001110100111101010010",
						 "101001110101001011110100",
						 "101001110101001010110110",
						 "101001110101001001111000",
						 "101001110101001000111010",
						 "101001110101000111111100",
						 "101001110101000110111110",
						 "101001110101000110000000",
						 "101001110101000101000010",
						 "101001110101000100000100",
						 "101001110101000011000110",
						 "101001110101000010001000",
						 "101001110101000001001010",
						 "101001110101000000001100",
						 "101001110100111111001110",
						 "101001110100111110010000",
						 "101001110100111101010010",
						 "101001110101001100000011",
						 "101001110101001011000100",
						 "101001110101001010000101",
						 "101001110101001001000110",
						 "101001110101001000000111",
						 "101001110101000111001000",
						 "101001110101000110001001",
						 "101001110101000101001010",
						 "101001110101000100001011",
						 "101001110101000011001100",
						 "101001110101000010001101",
						 "101001110101000001001110",
						 "101001110101000000001111",
						 "101001110100111111010000",
						 "101001110100111110010001",
						 "101001110100111101010010",
						 "101001110101001100000011",
						 "101001110101001011000100",
						 "101001110101001010000101",
						 "101001110101001001000110",
						 "101001110101001000000111",
						 "101001110101000111001000",
						 "101001110101000110001001",
						 "101001110101000101001010",
						 "101001110101000100001011",
						 "101001110101000011001100",
						 "101001110101000010001101",
						 "101001110101000001001110",
						 "101001110101000000001111",
						 "101001110100111111010000",
						 "101001110100111110010001",
						 "101001110100111101010010",
						 "101001110101001100000011",
						 "101001110101001011000100",
						 "101001110101001010000101",
						 "101001110101001001000110",
						 "101001110101001000000111",
						 "101001110101000111001000",
						 "101001110101000110001001",
						 "101001110101000101001010",
						 "101001110101000100001011",
						 "101001110101000011001100",
						 "101001110101000010001101",
						 "101001110101000001001110",
						 "101001110101000000001111",
						 "101001110100111111010000",
						 "101001110100111110010001",
						 "101001110100111101010010",
						 "101001110101001100010010",
						 "101001110101001011010010",
						 "101001110101001010010010",
						 "101001110101001001010010",
						 "101001110101001000010010",
						 "101001110101000111010010",
						 "101001110101000110010010",
						 "101001110101000101010010",
						 "101001110101000100010010",
						 "101001110101000011010010",
						 "101001110101000010010010",
						 "101001110101000001010010",
						 "101001110101000000010010",
						 "101001110100111111010010",
						 "101001110100111110010010",
						 "101001110100111101010010",
						 "101001110101001100010010",
						 "101001110101001011010010",
						 "101001110101001010010010",
						 "101001110101001001010010",
						 "101001110101001000010010",
						 "101001110101000111010010",
						 "101001110101000110010010",
						 "101001110101000101010010",
						 "101001110101000100010010",
						 "101001110101000011010010",
						 "101001110101000010010010",
						 "101001110101000001010010",
						 "101001110101000000010010",
						 "101001110100111111010010",
						 "101001110100111110010010",
						 "101001110100111101010010",
						 "101001110101001100010010",
						 "101001110101001011010010",
						 "101001110101001010010010",
						 "101001110101001001010010",
						 "101001110101001000010010",
						 "101001110101000111010010",
						 "101001110101000110010010",
						 "101001110101000101010010",
						 "101001110101000100010010",
						 "101001110101000011010010",
						 "101001110101000010010010",
						 "101001110101000001010010",
						 "101001110101000000010010",
						 "101001110100111111010010",
						 "101001110100111110010010",
						 "101001110100111101010010",
						 "101001110101001100100001",
						 "101001110101001011100000",
						 "101001110101001010011111",
						 "101001110101001001011110",
						 "101001110101001000011101",
						 "101001110101000111011100",
						 "101001110101000110011011",
						 "101001110101000101011010",
						 "101001110101000100011001",
						 "101001110101000011011000",
						 "101001110101000010010111",
						 "101001110101000001010110",
						 "101001110101000000010101",
						 "101001110100111111010100",
						 "101001110100111110010011",
						 "101001110100111101010010",
						 "101001110010101001100011",
						 "101001110010101000100010",
						 "101001110010100111100001",
						 "101001110010100110100000",
						 "101001110010100101011111",
						 "101001110010100100011110",
						 "101001110010100011011101",
						 "101001110010100010011100",
						 "101001110010100001011011",
						 "101001110010100000011010",
						 "101001110010011111011001",
						 "101001110010011110011000",
						 "101001110010011101010111",
						 "101001110010011100010110",
						 "101001110010011011010101",
						 "101001110010011010010100",
						 "101001110010101001110010",
						 "101001110010101000110000",
						 "101001110010100111101110",
						 "101001110010100110101100",
						 "101001110010100101101010",
						 "101001110010100100101000",
						 "101001110010100011100110",
						 "101001110010100010100100",
						 "101001110010100001100010",
						 "101001110010100000100000",
						 "101001110010011111011110",
						 "101001110010011110011100",
						 "101001110010011101011010",
						 "101001110010011100011000",
						 "101001110010011011010110",
						 "101001110010011010010100",
						 "101001110010101001110010",
						 "101001110010101000110000",
						 "101001110010100111101110",
						 "101001110010100110101100",
						 "101001110010100101101010",
						 "101001110010100100101000",
						 "101001110010100011100110",
						 "101001110010100010100100",
						 "101001110010100001100010",
						 "101001110010100000100000",
						 "101001110010011111011110",
						 "101001110010011110011100",
						 "101001110010011101011010",
						 "101001110010011100011000",
						 "101001110010011011010110",
						 "101001110010011010010100",
						 "101001110010101001110010",
						 "101001110010101000110000",
						 "101001110010100111101110",
						 "101001110010100110101100",
						 "101001110010100101101010",
						 "101001110010100100101000",
						 "101001110010100011100110",
						 "101001110010100010100100",
						 "101001110010100001100010",
						 "101001110010100000100000",
						 "101001110010011111011110",
						 "101001110010011110011100",
						 "101001110010011101011010",
						 "101001110010011100011000",
						 "101001110010011011010110",
						 "101001110010011010010100",
						 "101001110010101010000001",
						 "101001110010101000111110",
						 "101001110010100111111011",
						 "101001110010100110111000",
						 "101001110010100101110101",
						 "101001110010100100110010",
						 "101001110010100011101111",
						 "101001110010100010101100",
						 "101001110010100001101001",
						 "101001110010100000100110",
						 "101001110010011111100011",
						 "101001110010011110100000",
						 "101001110010011101011101",
						 "101001110010011100011010",
						 "101001110010011011010111",
						 "101001110010011010010100",
						 "101001110010101010000001",
						 "101001110010101000111110",
						 "101001110010100111111011",
						 "101001110010100110111000",
						 "101001110010100101110101",
						 "101001110010100100110010",
						 "101001110010100011101111",
						 "101001110010100010101100",
						 "101001110010100001101001",
						 "101001110010100000100110",
						 "101001110010011111100011",
						 "101001110010011110100000",
						 "101001110010011101011101",
						 "101001110010011100011010",
						 "101001110010011011010111",
						 "101001110010011010010100",
						 "101001110010101010000001",
						 "101001110010101000111110",
						 "101001110010100111111011",
						 "101001110010100110111000",
						 "101001110010100101110101",
						 "101001110010100100110010",
						 "101001110010100011101111",
						 "101001110010100010101100",
						 "101001110010100001101001",
						 "101001110010100000100110",
						 "101001110010011111100011",
						 "101001110010011110100000",
						 "101001110010011101011101",
						 "101001110010011100011010",
						 "101001110010011011010111",
						 "101001110010011010010100",
						 "101001110010101010010000",
						 "101001110010101001001100",
						 "101001110010101000001000",
						 "101001110010100111000100",
						 "101001110010100110000000",
						 "101001110010100100111100",
						 "101001110010100011111000",
						 "101001110010100010110100",
						 "101001110010100001110000",
						 "101001110010100000101100",
						 "101001110010011111101000",
						 "101001110010011110100100",
						 "101001110010011101100000",
						 "101001110010011100011100",
						 "101001110010011011011000",
						 "101001110010011010010100",
						 "101001110010101010010000",
						 "101001110010101001001100",
						 "101001110010101000001000",
						 "101001110010100111000100",
						 "101001110010100110000000",
						 "101001110010100100111100",
						 "101001110010100011111000",
						 "101001110010100010110100",
						 "101001110010100001110000",
						 "101001110010100000101100",
						 "101001110010011111101000",
						 "101001110010011110100100",
						 "101001110010011101100000",
						 "101001110010011100011100",
						 "101001110010011011011000",
						 "101001110010011010010100",
						 "101001110010101010011111",
						 "101001110010101001011010",
						 "101001110010101000010101",
						 "101001110010100111010000",
						 "101001110010100110001011",
						 "101001110010100101000110",
						 "101001110010100100000001",
						 "101001110010100010111100",
						 "101001110010100001110111",
						 "101001110010100000110010",
						 "101001110010011111101101",
						 "101001110010011110101000",
						 "101001110010011101100011",
						 "101001110010011100011110",
						 "101001110010011011011001",
						 "101001110010011010010100",
						 "101001110000000111100001",
						 "101001110000000110011100",
						 "101001110000000101010111",
						 "101001110000000100010010",
						 "101001110000000011001101",
						 "101001110000000010001000",
						 "101001110000000001000011",
						 "101001101111111111111110",
						 "101001101111111110111001",
						 "101001101111111101110100",
						 "101001101111111100101111",
						 "101001101111111011101010",
						 "101001101111111010100101",
						 "101001101111111001100000",
						 "101001101111111000011011",
						 "101001101111110111010110",
						 "101001110000000111100001",
						 "101001110000000110011100",
						 "101001110000000101010111",
						 "101001110000000100010010",
						 "101001110000000011001101",
						 "101001110000000010001000",
						 "101001110000000001000011",
						 "101001101111111111111110",
						 "101001101111111110111001",
						 "101001101111111101110100",
						 "101001101111111100101111",
						 "101001101111111011101010",
						 "101001101111111010100101",
						 "101001101111111001100000",
						 "101001101111111000011011",
						 "101001101111110111010110",
						 "101001110000000111110000",
						 "101001110000000110101010",
						 "101001110000000101100100",
						 "101001110000000100011110",
						 "101001110000000011011000",
						 "101001110000000010010010",
						 "101001110000000001001100",
						 "101001110000000000000110",
						 "101001101111111111000000",
						 "101001101111111101111010",
						 "101001101111111100110100",
						 "101001101111111011101110",
						 "101001101111111010101000",
						 "101001101111111001100010",
						 "101001101111111000011100",
						 "101001101111110111010110",
						 "101001110000000111110000",
						 "101001110000000110101010",
						 "101001110000000101100100",
						 "101001110000000100011110",
						 "101001110000000011011000",
						 "101001110000000010010010",
						 "101001110000000001001100",
						 "101001110000000000000110",
						 "101001101111111111000000",
						 "101001101111111101111010",
						 "101001101111111100110100",
						 "101001101111111011101110",
						 "101001101111111010101000",
						 "101001101111111001100010",
						 "101001101111111000011100",
						 "101001101111110111010110",
						 "101001110000000111110000",
						 "101001110000000110101010",
						 "101001110000000101100100",
						 "101001110000000100011110",
						 "101001110000000011011000",
						 "101001110000000010010010",
						 "101001110000000001001100",
						 "101001110000000000000110",
						 "101001101111111111000000",
						 "101001101111111101111010",
						 "101001101111111100110100",
						 "101001101111111011101110",
						 "101001101111111010101000",
						 "101001101111111001100010",
						 "101001101111111000011100",
						 "101001101111110111010110",
						 "101001110000000111111111",
						 "101001110000000110111000",
						 "101001110000000101110001",
						 "101001110000000100101010",
						 "101001110000000011100011",
						 "101001110000000010011100",
						 "101001110000000001010101",
						 "101001110000000000001110",
						 "101001101111111111000111",
						 "101001101111111110000000",
						 "101001101111111100111001",
						 "101001101111111011110010",
						 "101001101111111010101011",
						 "101001101111111001100100",
						 "101001101111111000011101",
						 "101001101111110111010110",
						 "101001110000000111111111",
						 "101001110000000110111000",
						 "101001110000000101110001",
						 "101001110000000100101010",
						 "101001110000000011100011",
						 "101001110000000010011100",
						 "101001110000000001010101",
						 "101001110000000000001110",
						 "101001101111111111000111",
						 "101001101111111110000000",
						 "101001101111111100111001",
						 "101001101111111011110010",
						 "101001101111111010101011",
						 "101001101111111001100100",
						 "101001101111111000011101",
						 "101001101111110111010110",
						 "101001110000001000001110",
						 "101001110000000111000110",
						 "101001110000000101111110",
						 "101001110000000100110110",
						 "101001110000000011101110",
						 "101001110000000010100110",
						 "101001110000000001011110",
						 "101001110000000000010110",
						 "101001101111111111001110",
						 "101001101111111110000110",
						 "101001101111111100111110",
						 "101001101111111011110110",
						 "101001101111111010101110",
						 "101001101111111001100110",
						 "101001101111111000011110",
						 "101001101111110111010110",
						 "101001110000001000001110",
						 "101001110000000111000110",
						 "101001110000000101111110",
						 "101001110000000100110110",
						 "101001110000000011101110",
						 "101001110000000010100110",
						 "101001110000000001011110",
						 "101001110000000000010110",
						 "101001101111111111001110",
						 "101001101111111110000110",
						 "101001101111111100111110",
						 "101001101111111011110110",
						 "101001101111111010101110",
						 "101001101111111001100110",
						 "101001101111111000011110",
						 "101001101111110111010110",
						 "101001101101100101010000",
						 "101001101101100100001000",
						 "101001101101100011000000",
						 "101001101101100001111000",
						 "101001101101100000110000",
						 "101001101101011111101000",
						 "101001101101011110100000",
						 "101001101101011101011000",
						 "101001101101011100010000",
						 "101001101101011011001000",
						 "101001101101011010000000",
						 "101001101101011000111000",
						 "101001101101010111110000",
						 "101001101101010110101000",
						 "101001101101010101100000",
						 "101001101101010100011000",
						 "101001101101100101011111",
						 "101001101101100100010110",
						 "101001101101100011001101",
						 "101001101101100010000100",
						 "101001101101100000111011",
						 "101001101101011111110010",
						 "101001101101011110101001",
						 "101001101101011101100000",
						 "101001101101011100010111",
						 "101001101101011011001110",
						 "101001101101011010000101",
						 "101001101101011000111100",
						 "101001101101010111110011",
						 "101001101101010110101010",
						 "101001101101010101100001",
						 "101001101101010100011000",
						 "101001101101100101011111",
						 "101001101101100100010110",
						 "101001101101100011001101",
						 "101001101101100010000100",
						 "101001101101100000111011",
						 "101001101101011111110010",
						 "101001101101011110101001",
						 "101001101101011101100000",
						 "101001101101011100010111",
						 "101001101101011011001110",
						 "101001101101011010000101",
						 "101001101101011000111100",
						 "101001101101010111110011",
						 "101001101101010110101010",
						 "101001101101010101100001",
						 "101001101101010100011000",
						 "101001101101100101011111",
						 "101001101101100100010110",
						 "101001101101100011001101",
						 "101001101101100010000100",
						 "101001101101100000111011",
						 "101001101101011111110010",
						 "101001101101011110101001",
						 "101001101101011101100000",
						 "101001101101011100010111",
						 "101001101101011011001110",
						 "101001101101011010000101",
						 "101001101101011000111100",
						 "101001101101010111110011",
						 "101001101101010110101010",
						 "101001101101010101100001",
						 "101001101101010100011000",
						 "101001101101100101101110",
						 "101001101101100100100100",
						 "101001101101100011011010",
						 "101001101101100010010000",
						 "101001101101100001000110",
						 "101001101101011111111100",
						 "101001101101011110110010",
						 "101001101101011101101000",
						 "101001101101011100011110",
						 "101001101101011011010100",
						 "101001101101011010001010",
						 "101001101101011001000000",
						 "101001101101010111110110",
						 "101001101101010110101100",
						 "101001101101010101100010",
						 "101001101101010100011000",
						 "101001101101100101101110",
						 "101001101101100100100100",
						 "101001101101100011011010",
						 "101001101101100010010000",
						 "101001101101100001000110",
						 "101001101101011111111100",
						 "101001101101011110110010",
						 "101001101101011101101000",
						 "101001101101011100011110",
						 "101001101101011011010100",
						 "101001101101011010001010",
						 "101001101101011001000000",
						 "101001101101010111110110",
						 "101001101101010110101100",
						 "101001101101010101100010",
						 "101001101101010100011000",
						 "101001101101100101111101",
						 "101001101101100100110010",
						 "101001101101100011100111",
						 "101001101101100010011100",
						 "101001101101100001010001",
						 "101001101101100000000110",
						 "101001101101011110111011",
						 "101001101101011101110000",
						 "101001101101011100100101",
						 "101001101101011011011010",
						 "101001101101011010001111",
						 "101001101101011001000100",
						 "101001101101010111111001",
						 "101001101101010110101110",
						 "101001101101010101100011",
						 "101001101101010100011000",
						 "101001101101100101111101",
						 "101001101101100100110010",
						 "101001101101100011100111",
						 "101001101101100010011100",
						 "101001101101100001010001",
						 "101001101101100000000110",
						 "101001101101011110111011",
						 "101001101101011101110000",
						 "101001101101011100100101",
						 "101001101101011011011010",
						 "101001101101011010001111",
						 "101001101101011001000100",
						 "101001101101010111111001",
						 "101001101101010110101110",
						 "101001101101010101100011",
						 "101001101101010100011000",
						 "101001101101100101111101",
						 "101001101101100100110010",
						 "101001101101100011100111",
						 "101001101101100010011100",
						 "101001101101100001010001",
						 "101001101101100000000110",
						 "101001101101011110111011",
						 "101001101101011101110000",
						 "101001101101011100100101",
						 "101001101101011011011010",
						 "101001101101011010001111",
						 "101001101101011001000100",
						 "101001101101010111111001",
						 "101001101101010110101110",
						 "101001101101010101100011",
						 "101001101101010100011000",
						 "101001101011000011001110",
						 "101001101011000010000010",
						 "101001101011000000110110",
						 "101001101010111111101010",
						 "101001101010111110011110",
						 "101001101010111101010010",
						 "101001101010111100000110",
						 "101001101010111010111010",
						 "101001101010111001101110",
						 "101001101010111000100010",
						 "101001101010110111010110",
						 "101001101010110110001010",
						 "101001101010110100111110",
						 "101001101010110011110010",
						 "101001101010110010100110",
						 "101001101010110001011010",
						 "101001101011000011001110",
						 "101001101011000010000010",
						 "101001101011000000110110",
						 "101001101010111111101010",
						 "101001101010111110011110",
						 "101001101010111101010010",
						 "101001101010111100000110",
						 "101001101010111010111010",
						 "101001101010111001101110",
						 "101001101010111000100010",
						 "101001101010110111010110",
						 "101001101010110110001010",
						 "101001101010110100111110",
						 "101001101010110011110010",
						 "101001101010110010100110",
						 "101001101010110001011010",
						 "101001101011000011001110",
						 "101001101011000010000010",
						 "101001101011000000110110",
						 "101001101010111111101010",
						 "101001101010111110011110",
						 "101001101010111101010010",
						 "101001101010111100000110",
						 "101001101010111010111010",
						 "101001101010111001101110",
						 "101001101010111000100010",
						 "101001101010110111010110",
						 "101001101010110110001010",
						 "101001101010110100111110",
						 "101001101010110011110010",
						 "101001101010110010100110",
						 "101001101010110001011010",
						 "101001101011000011011101",
						 "101001101011000010010000",
						 "101001101011000001000011",
						 "101001101010111111110110",
						 "101001101010111110101001",
						 "101001101010111101011100",
						 "101001101010111100001111",
						 "101001101010111011000010",
						 "101001101010111001110101",
						 "101001101010111000101000",
						 "101001101010110111011011",
						 "101001101010110110001110",
						 "101001101010110101000001",
						 "101001101010110011110100",
						 "101001101010110010100111",
						 "101001101010110001011010",
						 "101001101011000011011101",
						 "101001101011000010010000",
						 "101001101011000001000011",
						 "101001101010111111110110",
						 "101001101010111110101001",
						 "101001101010111101011100",
						 "101001101010111100001111",
						 "101001101010111011000010",
						 "101001101010111001110101",
						 "101001101010111000101000",
						 "101001101010110111011011",
						 "101001101010110110001110",
						 "101001101010110101000001",
						 "101001101010110011110100",
						 "101001101010110010100111",
						 "101001101010110001011010",
						 "101001101011000011101100",
						 "101001101011000010011110",
						 "101001101011000001010000",
						 "101001101011000000000010",
						 "101001101010111110110100",
						 "101001101010111101100110",
						 "101001101010111100011000",
						 "101001101010111011001010",
						 "101001101010111001111100",
						 "101001101010111000101110",
						 "101001101010110111100000",
						 "101001101010110110010010",
						 "101001101010110101000100",
						 "101001101010110011110110",
						 "101001101010110010101000",
						 "101001101010110001011010",
						 "101001101011000011101100",
						 "101001101011000010011110",
						 "101001101011000001010000",
						 "101001101011000000000010",
						 "101001101010111110110100",
						 "101001101010111101100110",
						 "101001101010111100011000",
						 "101001101010111011001010",
						 "101001101010111001111100",
						 "101001101010111000101110",
						 "101001101010110111100000",
						 "101001101010110110010010",
						 "101001101010110101000100",
						 "101001101010110011110110",
						 "101001101010110010101000",
						 "101001101010110001011010",
						 "101001101011000011101100",
						 "101001101011000010011110",
						 "101001101011000001010000",
						 "101001101011000000000010",
						 "101001101010111110110100",
						 "101001101010111101100110",
						 "101001101010111100011000",
						 "101001101010111011001010",
						 "101001101010111001111100",
						 "101001101010111000101110",
						 "101001101010110111100000",
						 "101001101010110110010010",
						 "101001101010110101000100",
						 "101001101010110011110110",
						 "101001101010110010101000",
						 "101001101010110001011010",
						 "101001101000100000111101",
						 "101001101000011111101110",
						 "101001101000011110011111",
						 "101001101000011101010000",
						 "101001101000011100000001",
						 "101001101000011010110010",
						 "101001101000011001100011",
						 "101001101000011000010100",
						 "101001101000010111000101",
						 "101001101000010101110110",
						 "101001101000010100100111",
						 "101001101000010011011000",
						 "101001101000010010001001",
						 "101001101000010000111010",
						 "101001101000001111101011",
						 "101001101000001110011100",
						 "101001101000100000111101",
						 "101001101000011111101110",
						 "101001101000011110011111",
						 "101001101000011101010000",
						 "101001101000011100000001",
						 "101001101000011010110010",
						 "101001101000011001100011",
						 "101001101000011000010100",
						 "101001101000010111000101",
						 "101001101000010101110110",
						 "101001101000010100100111",
						 "101001101000010011011000",
						 "101001101000010010001001",
						 "101001101000010000111010",
						 "101001101000001111101011",
						 "101001101000001110011100",
						 "101001101000100000111101",
						 "101001101000011111101110",
						 "101001101000011110011111",
						 "101001101000011101010000",
						 "101001101000011100000001",
						 "101001101000011010110010",
						 "101001101000011001100011",
						 "101001101000011000010100",
						 "101001101000010111000101",
						 "101001101000010101110110",
						 "101001101000010100100111",
						 "101001101000010011011000",
						 "101001101000010010001001",
						 "101001101000010000111010",
						 "101001101000001111101011",
						 "101001101000001110011100",
						 "101001101000100001001100",
						 "101001101000011111111100",
						 "101001101000011110101100",
						 "101001101000011101011100",
						 "101001101000011100001100",
						 "101001101000011010111100",
						 "101001101000011001101100",
						 "101001101000011000011100",
						 "101001101000010111001100",
						 "101001101000010101111100",
						 "101001101000010100101100",
						 "101001101000010011011100",
						 "101001101000010010001100",
						 "101001101000010000111100",
						 "101001101000001111101100",
						 "101001101000001110011100",
						 "101001101000100001001100",
						 "101001101000011111111100",
						 "101001101000011110101100",
						 "101001101000011101011100",
						 "101001101000011100001100",
						 "101001101000011010111100",
						 "101001101000011001101100",
						 "101001101000011000011100",
						 "101001101000010111001100",
						 "101001101000010101111100",
						 "101001101000010100101100",
						 "101001101000010011011100",
						 "101001101000010010001100",
						 "101001101000010000111100",
						 "101001101000001111101100",
						 "101001101000001110011100",
						 "101001101000100001011011",
						 "101001101000100000001010",
						 "101001101000011110111001",
						 "101001101000011101101000",
						 "101001101000011100010111",
						 "101001101000011011000110",
						 "101001101000011001110101",
						 "101001101000011000100100",
						 "101001101000010111010011",
						 "101001101000010110000010",
						 "101001101000010100110001",
						 "101001101000010011100000",
						 "101001101000010010001111",
						 "101001101000010000111110",
						 "101001101000001111101101",
						 "101001101000001110011100",
						 "101001101000100001011011",
						 "101001101000100000001010",
						 "101001101000011110111001",
						 "101001101000011101101000",
						 "101001101000011100010111",
						 "101001101000011011000110",
						 "101001101000011001110101",
						 "101001101000011000100100",
						 "101001101000010111010011",
						 "101001101000010110000010",
						 "101001101000010100110001",
						 "101001101000010011100000",
						 "101001101000010010001111",
						 "101001101000010000111110",
						 "101001101000001111101101",
						 "101001101000001110011100",
						 "101001101000100001011011",
						 "101001101000100000001010",
						 "101001101000011110111001",
						 "101001101000011101101000",
						 "101001101000011100010111",
						 "101001101000011011000110",
						 "101001101000011001110101",
						 "101001101000011000100100",
						 "101001101000010111010011",
						 "101001101000010110000010",
						 "101001101000010100110001",
						 "101001101000010011100000",
						 "101001101000010010001111",
						 "101001101000010000111110",
						 "101001101000001111101101",
						 "101001101000001110011100",
						 "101001101000100001101010",
						 "101001101000100000011000",
						 "101001101000011111000110",
						 "101001101000011101110100",
						 "101001101000011100100010",
						 "101001101000011011010000",
						 "101001101000011001111110",
						 "101001101000011000101100",
						 "101001101000010111011010",
						 "101001101000010110001000",
						 "101001101000010100110110",
						 "101001101000010011100100",
						 "101001101000010010010010",
						 "101001101000010001000000",
						 "101001101000001111101110",
						 "101001101000001110011100",
						 "101001100101111110101100",
						 "101001100101111101011010",
						 "101001100101111100001000",
						 "101001100101111010110110",
						 "101001100101111001100100",
						 "101001100101111000010010",
						 "101001100101110111000000",
						 "101001100101110101101110",
						 "101001100101110100011100",
						 "101001100101110011001010",
						 "101001100101110001111000",
						 "101001100101110000100110",
						 "101001100101101111010100",
						 "101001100101101110000010",
						 "101001100101101100110000",
						 "101001100101101011011110",
						 "101001100101111110101100",
						 "101001100101111101011010",
						 "101001100101111100001000",
						 "101001100101111010110110",
						 "101001100101111001100100",
						 "101001100101111000010010",
						 "101001100101110111000000",
						 "101001100101110101101110",
						 "101001100101110100011100",
						 "101001100101110011001010",
						 "101001100101110001111000",
						 "101001100101110000100110",
						 "101001100101101111010100",
						 "101001100101101110000010",
						 "101001100101101100110000",
						 "101001100101101011011110",
						 "101001100101111110111011",
						 "101001100101111101101000",
						 "101001100101111100010101",
						 "101001100101111011000010",
						 "101001100101111001101111",
						 "101001100101111000011100",
						 "101001100101110111001001",
						 "101001100101110101110110",
						 "101001100101110100100011",
						 "101001100101110011010000",
						 "101001100101110001111101",
						 "101001100101110000101010",
						 "101001100101101111010111",
						 "101001100101101110000100",
						 "101001100101101100110001",
						 "101001100101101011011110",
						 "101001100101111110111011",
						 "101001100101111101101000",
						 "101001100101111100010101",
						 "101001100101111011000010",
						 "101001100101111001101111",
						 "101001100101111000011100",
						 "101001100101110111001001",
						 "101001100101110101110110",
						 "101001100101110100100011",
						 "101001100101110011010000",
						 "101001100101110001111101",
						 "101001100101110000101010",
						 "101001100101101111010111",
						 "101001100101101110000100",
						 "101001100101101100110001",
						 "101001100101101011011110",
						 "101001100101111110111011",
						 "101001100101111101101000",
						 "101001100101111100010101",
						 "101001100101111011000010",
						 "101001100101111001101111",
						 "101001100101111000011100",
						 "101001100101110111001001",
						 "101001100101110101110110",
						 "101001100101110100100011",
						 "101001100101110011010000",
						 "101001100101110001111101",
						 "101001100101110000101010",
						 "101001100101101111010111",
						 "101001100101101110000100",
						 "101001100101101100110001",
						 "101001100101101011011110",
						 "101001100101111111001010",
						 "101001100101111101110110",
						 "101001100101111100100010",
						 "101001100101111011001110",
						 "101001100101111001111010",
						 "101001100101111000100110",
						 "101001100101110111010010",
						 "101001100101110101111110",
						 "101001100101110100101010",
						 "101001100101110011010110",
						 "101001100101110010000010",
						 "101001100101110000101110",
						 "101001100101101111011010",
						 "101001100101101110000110",
						 "101001100101101100110010",
						 "101001100101101011011110",
						 "101001100101111111001010",
						 "101001100101111101110110",
						 "101001100101111100100010",
						 "101001100101111011001110",
						 "101001100101111001111010",
						 "101001100101111000100110",
						 "101001100101110111010010",
						 "101001100101110101111110",
						 "101001100101110100101010",
						 "101001100101110011010110",
						 "101001100101110010000010",
						 "101001100101110000101110",
						 "101001100101101111011010",
						 "101001100101101110000110",
						 "101001100101101100110010",
						 "101001100101101011011110",
						 "101001100011011100011011",
						 "101001100011011011000110",
						 "101001100011011001110001",
						 "101001100011011000011100",
						 "101001100011010111000111",
						 "101001100011010101110010",
						 "101001100011010100011101",
						 "101001100011010011001000",
						 "101001100011010001110011",
						 "101001100011010000011110",
						 "101001100011001111001001",
						 "101001100011001101110100",
						 "101001100011001100011111",
						 "101001100011001011001010",
						 "101001100011001001110101",
						 "101001100011001000100000",
						 "101001100011011100011011",
						 "101001100011011011000110",
						 "101001100011011001110001",
						 "101001100011011000011100",
						 "101001100011010111000111",
						 "101001100011010101110010",
						 "101001100011010100011101",
						 "101001100011010011001000",
						 "101001100011010001110011",
						 "101001100011010000011110",
						 "101001100011001111001001",
						 "101001100011001101110100",
						 "101001100011001100011111",
						 "101001100011001011001010",
						 "101001100011001001110101",
						 "101001100011001000100000",
						 "101001100011011100011011",
						 "101001100011011011000110",
						 "101001100011011001110001",
						 "101001100011011000011100",
						 "101001100011010111000111",
						 "101001100011010101110010",
						 "101001100011010100011101",
						 "101001100011010011001000",
						 "101001100011010001110011",
						 "101001100011010000011110",
						 "101001100011001111001001",
						 "101001100011001101110100",
						 "101001100011001100011111",
						 "101001100011001011001010",
						 "101001100011001001110101",
						 "101001100011001000100000",
						 "101001100011011100101010",
						 "101001100011011011010100",
						 "101001100011011001111110",
						 "101001100011011000101000",
						 "101001100011010111010010",
						 "101001100011010101111100",
						 "101001100011010100100110",
						 "101001100011010011010000",
						 "101001100011010001111010",
						 "101001100011010000100100",
						 "101001100011001111001110",
						 "101001100011001101111000",
						 "101001100011001100100010",
						 "101001100011001011001100",
						 "101001100011001001110110",
						 "101001100011001000100000",
						 "101001100011011100101010",
						 "101001100011011011010100",
						 "101001100011011001111110",
						 "101001100011011000101000",
						 "101001100011010111010010",
						 "101001100011010101111100",
						 "101001100011010100100110",
						 "101001100011010011010000",
						 "101001100011010001111010",
						 "101001100011010000100100",
						 "101001100011001111001110",
						 "101001100011001101111000",
						 "101001100011001100100010",
						 "101001100011001011001100",
						 "101001100011001001110110",
						 "101001100011001000100000",
						 "101001100011011100101010",
						 "101001100011011011010100",
						 "101001100011011001111110",
						 "101001100011011000101000",
						 "101001100011010111010010",
						 "101001100011010101111100",
						 "101001100011010100100110",
						 "101001100011010011010000",
						 "101001100011010001111010",
						 "101001100011010000100100",
						 "101001100011001111001110",
						 "101001100011001101111000",
						 "101001100011001100100010",
						 "101001100011001011001100",
						 "101001100011001001110110",
						 "101001100011001000100000",
						 "101001100011011100111001",
						 "101001100011011011100010",
						 "101001100011011010001011",
						 "101001100011011000110100",
						 "101001100011010111011101",
						 "101001100011010110000110",
						 "101001100011010100101111",
						 "101001100011010011011000",
						 "101001100011010010000001",
						 "101001100011010000101010",
						 "101001100011001111010011",
						 "101001100011001101111100",
						 "101001100011001100100101",
						 "101001100011001011001110",
						 "101001100011001001110111",
						 "101001100011001000100000",
						 "101001100011011100111001",
						 "101001100011011011100010",
						 "101001100011011010001011",
						 "101001100011011000110100",
						 "101001100011010111011101",
						 "101001100011010110000110",
						 "101001100011010100101111",
						 "101001100011010011011000",
						 "101001100011010010000001",
						 "101001100011010000101010",
						 "101001100011001111010011",
						 "101001100011001101111100",
						 "101001100011001100100101",
						 "101001100011001011001110",
						 "101001100011001001110111",
						 "101001100011001000100000",
						 "101001100000111010001010",
						 "101001100000111000110010",
						 "101001100000110111011010",
						 "101001100000110110000010",
						 "101001100000110100101010",
						 "101001100000110011010010",
						 "101001100000110001111010",
						 "101001100000110000100010",
						 "101001100000101111001010",
						 "101001100000101101110010",
						 "101001100000101100011010",
						 "101001100000101011000010",
						 "101001100000101001101010",
						 "101001100000101000010010",
						 "101001100000100110111010",
						 "101001100000100101100010",
						 "101001100000111010001010",
						 "101001100000111000110010",
						 "101001100000110111011010",
						 "101001100000110110000010",
						 "101001100000110100101010",
						 "101001100000110011010010",
						 "101001100000110001111010",
						 "101001100000110000100010",
						 "101001100000101111001010",
						 "101001100000101101110010",
						 "101001100000101100011010",
						 "101001100000101011000010",
						 "101001100000101001101010",
						 "101001100000101000010010",
						 "101001100000100110111010",
						 "101001100000100101100010",
						 "101001100000111010001010",
						 "101001100000111000110010",
						 "101001100000110111011010",
						 "101001100000110110000010",
						 "101001100000110100101010",
						 "101001100000110011010010",
						 "101001100000110001111010",
						 "101001100000110000100010",
						 "101001100000101111001010",
						 "101001100000101101110010",
						 "101001100000101100011010",
						 "101001100000101011000010",
						 "101001100000101001101010",
						 "101001100000101000010010",
						 "101001100000100110111010",
						 "101001100000100101100010",
						 "101001100000111010011001",
						 "101001100000111001000000",
						 "101001100000110111100111",
						 "101001100000110110001110",
						 "101001100000110100110101",
						 "101001100000110011011100",
						 "101001100000110010000011",
						 "101001100000110000101010",
						 "101001100000101111010001",
						 "101001100000101101111000",
						 "101001100000101100011111",
						 "101001100000101011000110",
						 "101001100000101001101101",
						 "101001100000101000010100",
						 "101001100000100110111011",
						 "101001100000100101100010",
						 "101001100000111010011001",
						 "101001100000111001000000",
						 "101001100000110111100111",
						 "101001100000110110001110",
						 "101001100000110100110101",
						 "101001100000110011011100",
						 "101001100000110010000011",
						 "101001100000110000101010",
						 "101001100000101111010001",
						 "101001100000101101111000",
						 "101001100000101100011111",
						 "101001100000101011000110",
						 "101001100000101001101101",
						 "101001100000101000010100",
						 "101001100000100110111011",
						 "101001100000100101100010",
						 "101001100000111010011001",
						 "101001100000111001000000",
						 "101001100000110111100111",
						 "101001100000110110001110",
						 "101001100000110100110101",
						 "101001100000110011011100",
						 "101001100000110010000011",
						 "101001100000110000101010",
						 "101001100000101111010001",
						 "101001100000101101111000",
						 "101001100000101100011111",
						 "101001100000101011000110",
						 "101001100000101001101101",
						 "101001100000101000010100",
						 "101001100000100110111011",
						 "101001100000100101100010",
						 "101001100000111010101000",
						 "101001100000111001001110",
						 "101001100000110111110100",
						 "101001100000110110011010",
						 "101001100000110101000000",
						 "101001100000110011100110",
						 "101001100000110010001100",
						 "101001100000110000110010",
						 "101001100000101111011000",
						 "101001100000101101111110",
						 "101001100000101100100100",
						 "101001100000101011001010",
						 "101001100000101001110000",
						 "101001100000101000010110",
						 "101001100000100110111100",
						 "101001100000100101100010",
						 "101001011110010111101010",
						 "101001011110010110010000",
						 "101001011110010100110110",
						 "101001011110010011011100",
						 "101001011110010010000010",
						 "101001011110010000101000",
						 "101001011110001111001110",
						 "101001011110001101110100",
						 "101001011110001100011010",
						 "101001011110001011000000",
						 "101001011110001001100110",
						 "101001011110001000001100",
						 "101001011110000110110010",
						 "101001011110000101011000",
						 "101001011110000011111110",
						 "101001011110000010100100",
						 "101001011110010111101010",
						 "101001011110010110010000",
						 "101001011110010100110110",
						 "101001011110010011011100",
						 "101001011110010010000010",
						 "101001011110010000101000",
						 "101001011110001111001110",
						 "101001011110001101110100",
						 "101001011110001100011010",
						 "101001011110001011000000",
						 "101001011110001001100110",
						 "101001011110001000001100",
						 "101001011110000110110010",
						 "101001011110000101011000",
						 "101001011110000011111110",
						 "101001011110000010100100",
						 "101001011110010111111001",
						 "101001011110010110011110",
						 "101001011110010101000011",
						 "101001011110010011101000",
						 "101001011110010010001101",
						 "101001011110010000110010",
						 "101001011110001111010111",
						 "101001011110001101111100",
						 "101001011110001100100001",
						 "101001011110001011000110",
						 "101001011110001001101011",
						 "101001011110001000010000",
						 "101001011110000110110101",
						 "101001011110000101011010",
						 "101001011110000011111111",
						 "101001011110000010100100",
						 "101001011110010111111001",
						 "101001011110010110011110",
						 "101001011110010101000011",
						 "101001011110010011101000",
						 "101001011110010010001101",
						 "101001011110010000110010",
						 "101001011110001111010111",
						 "101001011110001101111100",
						 "101001011110001100100001",
						 "101001011110001011000110",
						 "101001011110001001101011",
						 "101001011110001000010000",
						 "101001011110000110110101",
						 "101001011110000101011010",
						 "101001011110000011111111",
						 "101001011110000010100100",
						 "101001011110011000001000",
						 "101001011110010110101100",
						 "101001011110010101010000",
						 "101001011110010011110100",
						 "101001011110010010011000",
						 "101001011110010000111100",
						 "101001011110001111100000",
						 "101001011110001110000100",
						 "101001011110001100101000",
						 "101001011110001011001100",
						 "101001011110001001110000",
						 "101001011110001000010100",
						 "101001011110000110111000",
						 "101001011110000101011100",
						 "101001011110000100000000",
						 "101001011110000010100100",
						 "101001011110011000001000",
						 "101001011110010110101100",
						 "101001011110010101010000",
						 "101001011110010011110100",
						 "101001011110010010011000",
						 "101001011110010000111100",
						 "101001011110001111100000",
						 "101001011110001110000100",
						 "101001011110001100101000",
						 "101001011110001011001100",
						 "101001011110001001110000",
						 "101001011110001000010100",
						 "101001011110000110111000",
						 "101001011110000101011100",
						 "101001011110000100000000",
						 "101001011110000010100100",
						 "101001011110011000001000",
						 "101001011110010110101100",
						 "101001011110010101010000",
						 "101001011110010011110100",
						 "101001011110010010011000",
						 "101001011110010000111100",
						 "101001011110001111100000",
						 "101001011110001110000100",
						 "101001011110001100101000",
						 "101001011110001011001100",
						 "101001011110001001110000",
						 "101001011110001000010100",
						 "101001011110000110111000",
						 "101001011110000101011100",
						 "101001011110000100000000",
						 "101001011110000010100100",
						 "101001011011110101011001",
						 "101001011011110011111100",
						 "101001011011110010011111",
						 "101001011011110001000010",
						 "101001011011101111100101",
						 "101001011011101110001000",
						 "101001011011101100101011",
						 "101001011011101011001110",
						 "101001011011101001110001",
						 "101001011011101000010100",
						 "101001011011100110110111",
						 "101001011011100101011010",
						 "101001011011100011111101",
						 "101001011011100010100000",
						 "101001011011100001000011",
						 "101001011011011111100110",
						 "101001011011110101011001",
						 "101001011011110011111100",
						 "101001011011110010011111",
						 "101001011011110001000010",
						 "101001011011101111100101",
						 "101001011011101110001000",
						 "101001011011101100101011",
						 "101001011011101011001110",
						 "101001011011101001110001",
						 "101001011011101000010100",
						 "101001011011100110110111",
						 "101001011011100101011010",
						 "101001011011100011111101",
						 "101001011011100010100000",
						 "101001011011100001000011",
						 "101001011011011111100110",
						 "101001011011110101011001",
						 "101001011011110011111100",
						 "101001011011110010011111",
						 "101001011011110001000010",
						 "101001011011101111100101",
						 "101001011011101110001000",
						 "101001011011101100101011",
						 "101001011011101011001110",
						 "101001011011101001110001",
						 "101001011011101000010100",
						 "101001011011100110110111",
						 "101001011011100101011010",
						 "101001011011100011111101",
						 "101001011011100010100000",
						 "101001011011100001000011",
						 "101001011011011111100110",
						 "101001011011110101101000",
						 "101001011011110100001010",
						 "101001011011110010101100",
						 "101001011011110001001110",
						 "101001011011101111110000",
						 "101001011011101110010010",
						 "101001011011101100110100",
						 "101001011011101011010110",
						 "101001011011101001111000",
						 "101001011011101000011010",
						 "101001011011100110111100",
						 "101001011011100101011110",
						 "101001011011100100000000",
						 "101001011011100010100010",
						 "101001011011100001000100",
						 "101001011011011111100110",
						 "101001011011110101101000",
						 "101001011011110100001010",
						 "101001011011110010101100",
						 "101001011011110001001110",
						 "101001011011101111110000",
						 "101001011011101110010010",
						 "101001011011101100110100",
						 "101001011011101011010110",
						 "101001011011101001111000",
						 "101001011011101000011010",
						 "101001011011100110111100",
						 "101001011011100101011110",
						 "101001011011100100000000",
						 "101001011011100010100010",
						 "101001011011100001000100",
						 "101001011011011111100110",
						 "101001011011110101101000",
						 "101001011011110100001010",
						 "101001011011110010101100",
						 "101001011011110001001110",
						 "101001011011101111110000",
						 "101001011011101110010010",
						 "101001011011101100110100",
						 "101001011011101011010110",
						 "101001011011101001111000",
						 "101001011011101000011010",
						 "101001011011100110111100",
						 "101001011011100101011110",
						 "101001011011100100000000",
						 "101001011011100010100010",
						 "101001011011100001000100",
						 "101001011011011111100110",
						 "101001011011110101110111",
						 "101001011011110100011000",
						 "101001011011110010111001",
						 "101001011011110001011010",
						 "101001011011101111111011",
						 "101001011011101110011100",
						 "101001011011101100111101",
						 "101001011011101011011110",
						 "101001011011101001111111",
						 "101001011011101000100000",
						 "101001011011100111000001",
						 "101001011011100101100010",
						 "101001011011100100000011",
						 "101001011011100010100100",
						 "101001011011100001000101",
						 "101001011011011111100110",
						 "101001011001010010111001",
						 "101001011001010001011010",
						 "101001011001001111111011",
						 "101001011001001110011100",
						 "101001011001001100111101",
						 "101001011001001011011110",
						 "101001011001001001111111",
						 "101001011001001000100000",
						 "101001011001000111000001",
						 "101001011001000101100010",
						 "101001011001000100000011",
						 "101001011001000010100100",
						 "101001011001000001000101",
						 "101001011000111111100110",
						 "101001011000111110000111",
						 "101001011000111100101000",
						 "101001011001010011001000",
						 "101001011001010001101000",
						 "101001011001010000001000",
						 "101001011001001110101000",
						 "101001011001001101001000",
						 "101001011001001011101000",
						 "101001011001001010001000",
						 "101001011001001000101000",
						 "101001011001000111001000",
						 "101001011001000101101000",
						 "101001011001000100001000",
						 "101001011001000010101000",
						 "101001011001000001001000",
						 "101001011000111111101000",
						 "101001011000111110001000",
						 "101001011000111100101000",
						 "101001011001010011001000",
						 "101001011001010001101000",
						 "101001011001010000001000",
						 "101001011001001110101000",
						 "101001011001001101001000",
						 "101001011001001011101000",
						 "101001011001001010001000",
						 "101001011001001000101000",
						 "101001011001000111001000",
						 "101001011001000101101000",
						 "101001011001000100001000",
						 "101001011001000010101000",
						 "101001011001000001001000",
						 "101001011000111111101000",
						 "101001011000111110001000",
						 "101001011000111100101000",
						 "101001011001010011001000",
						 "101001011001010001101000",
						 "101001011001010000001000",
						 "101001011001001110101000",
						 "101001011001001101001000",
						 "101001011001001011101000",
						 "101001011001001010001000",
						 "101001011001001000101000",
						 "101001011001000111001000",
						 "101001011001000101101000",
						 "101001011001000100001000",
						 "101001011001000010101000",
						 "101001011001000001001000",
						 "101001011000111111101000",
						 "101001011000111110001000",
						 "101001011000111100101000",
						 "101001011001010011010111",
						 "101001011001010001110110",
						 "101001011001010000010101",
						 "101001011001001110110100",
						 "101001011001001101010011",
						 "101001011001001011110010",
						 "101001011001001010010001",
						 "101001011001001000110000",
						 "101001011001000111001111",
						 "101001011001000101101110",
						 "101001011001000100001101",
						 "101001011001000010101100",
						 "101001011001000001001011",
						 "101001011000111111101010",
						 "101001011000111110001001",
						 "101001011000111100101000",
						 "101001011001010011010111",
						 "101001011001010001110110",
						 "101001011001010000010101",
						 "101001011001001110110100",
						 "101001011001001101010011",
						 "101001011001001011110010",
						 "101001011001001010010001",
						 "101001011001001000110000",
						 "101001011001000111001111",
						 "101001011001000101101110",
						 "101001011001000100001101",
						 "101001011001000010101100",
						 "101001011001000001001011",
						 "101001011000111111101010",
						 "101001011000111110001001",
						 "101001011000111100101000",
						 "101001011001010011010111",
						 "101001011001010001110110",
						 "101001011001010000010101",
						 "101001011001001110110100",
						 "101001011001001101010011",
						 "101001011001001011110010",
						 "101001011001001010010001",
						 "101001011001001000110000",
						 "101001011001000111001111",
						 "101001011001000101101110",
						 "101001011001000100001101",
						 "101001011001000010101100",
						 "101001011001000001001011",
						 "101001011000111111101010",
						 "101001011000111110001001",
						 "101001011000111100101000",
						 "101001010110110000101000",
						 "101001010110101111000110",
						 "101001010110101101100100",
						 "101001010110101100000010",
						 "101001010110101010100000",
						 "101001010110101000111110",
						 "101001010110100111011100",
						 "101001010110100101111010",
						 "101001010110100100011000",
						 "101001010110100010110110",
						 "101001010110100001010100",
						 "101001010110011111110010",
						 "101001010110011110010000",
						 "101001010110011100101110",
						 "101001010110011011001100",
						 "101001010110011001101010",
						 "101001010110110000101000",
						 "101001010110101111000110",
						 "101001010110101101100100",
						 "101001010110101100000010",
						 "101001010110101010100000",
						 "101001010110101000111110",
						 "101001010110100111011100",
						 "101001010110100101111010",
						 "101001010110100100011000",
						 "101001010110100010110110",
						 "101001010110100001010100",
						 "101001010110011111110010",
						 "101001010110011110010000",
						 "101001010110011100101110",
						 "101001010110011011001100",
						 "101001010110011001101010",
						 "101001010110110000101000",
						 "101001010110101111000110",
						 "101001010110101101100100",
						 "101001010110101100000010",
						 "101001010110101010100000",
						 "101001010110101000111110",
						 "101001010110100111011100",
						 "101001010110100101111010",
						 "101001010110100100011000",
						 "101001010110100010110110",
						 "101001010110100001010100",
						 "101001010110011111110010",
						 "101001010110011110010000",
						 "101001010110011100101110",
						 "101001010110011011001100",
						 "101001010110011001101010",
						 "101001010110110000110111",
						 "101001010110101111010100",
						 "101001010110101101110001",
						 "101001010110101100001110",
						 "101001010110101010101011",
						 "101001010110101001001000",
						 "101001010110100111100101",
						 "101001010110100110000010",
						 "101001010110100100011111",
						 "101001010110100010111100",
						 "101001010110100001011001",
						 "101001010110011111110110",
						 "101001010110011110010011",
						 "101001010110011100110000",
						 "101001010110011011001101",
						 "101001010110011001101010",
						 "101001010110110000110111",
						 "101001010110101111010100",
						 "101001010110101101110001",
						 "101001010110101100001110",
						 "101001010110101010101011",
						 "101001010110101001001000",
						 "101001010110100111100101",
						 "101001010110100110000010",
						 "101001010110100100011111",
						 "101001010110100010111100",
						 "101001010110100001011001",
						 "101001010110011111110110",
						 "101001010110011110010011",
						 "101001010110011100110000",
						 "101001010110011011001101",
						 "101001010110011001101010",
						 "101001010110110001000110",
						 "101001010110101111100010",
						 "101001010110101101111110",
						 "101001010110101100011010",
						 "101001010110101010110110",
						 "101001010110101001010010",
						 "101001010110100111101110",
						 "101001010110100110001010",
						 "101001010110100100100110",
						 "101001010110100011000010",
						 "101001010110100001011110",
						 "101001010110011111111010",
						 "101001010110011110010110",
						 "101001010110011100110010",
						 "101001010110011011001110",
						 "101001010110011001101010",
						 "101001010110110001000110",
						 "101001010110101111100010",
						 "101001010110101101111110",
						 "101001010110101100011010",
						 "101001010110101010110110",
						 "101001010110101001010010",
						 "101001010110100111101110",
						 "101001010110100110001010",
						 "101001010110100100100110",
						 "101001010110100011000010",
						 "101001010110100001011110",
						 "101001010110011111111010",
						 "101001010110011110010110",
						 "101001010110011100110010",
						 "101001010110011011001110",
						 "101001010110011001101010",
						 "101001010100001110001000",
						 "101001010100001100100100",
						 "101001010100001011000000",
						 "101001010100001001011100",
						 "101001010100000111111000",
						 "101001010100000110010100",
						 "101001010100000100110000",
						 "101001010100000011001100",
						 "101001010100000001101000",
						 "101001010100000000000100",
						 "101001010011111110100000",
						 "101001010011111100111100",
						 "101001010011111011011000",
						 "101001010011111001110100",
						 "101001010011111000010000",
						 "101001010011110110101100",
						 "101001010100001110010111",
						 "101001010100001100110010",
						 "101001010100001011001101",
						 "101001010100001001101000",
						 "101001010100001000000011",
						 "101001010100000110011110",
						 "101001010100000100111001",
						 "101001010100000011010100",
						 "101001010100000001101111",
						 "101001010100000000001010",
						 "101001010011111110100101",
						 "101001010011111101000000",
						 "101001010011111011011011",
						 "101001010011111001110110",
						 "101001010011111000010001",
						 "101001010011110110101100",
						 "101001010100001110010111",
						 "101001010100001100110010",
						 "101001010100001011001101",
						 "101001010100001001101000",
						 "101001010100001000000011",
						 "101001010100000110011110",
						 "101001010100000100111001",
						 "101001010100000011010100",
						 "101001010100000001101111",
						 "101001010100000000001010",
						 "101001010011111110100101",
						 "101001010011111101000000",
						 "101001010011111011011011",
						 "101001010011111001110110",
						 "101001010011111000010001",
						 "101001010011110110101100",
						 "101001010100001110010111",
						 "101001010100001100110010",
						 "101001010100001011001101",
						 "101001010100001001101000",
						 "101001010100001000000011",
						 "101001010100000110011110",
						 "101001010100000100111001",
						 "101001010100000011010100",
						 "101001010100000001101111",
						 "101001010100000000001010",
						 "101001010011111110100101",
						 "101001010011111101000000",
						 "101001010011111011011011",
						 "101001010011111001110110",
						 "101001010011111000010001",
						 "101001010011110110101100",
						 "101001010100001110100110",
						 "101001010100001101000000",
						 "101001010100001011011010",
						 "101001010100001001110100",
						 "101001010100001000001110",
						 "101001010100000110101000",
						 "101001010100000101000010",
						 "101001010100000011011100",
						 "101001010100000001110110",
						 "101001010100000000010000",
						 "101001010011111110101010",
						 "101001010011111101000100",
						 "101001010011111011011110",
						 "101001010011111001111000",
						 "101001010011111000010010",
						 "101001010011110110101100",
						 "101001010100001110100110",
						 "101001010100001101000000",
						 "101001010100001011011010",
						 "101001010100001001110100",
						 "101001010100001000001110",
						 "101001010100000110101000",
						 "101001010100000101000010",
						 "101001010100000011011100",
						 "101001010100000001110110",
						 "101001010100000000010000",
						 "101001010011111110101010",
						 "101001010011111101000100",
						 "101001010011111011011110",
						 "101001010011111001111000",
						 "101001010011111000010010",
						 "101001010011110110101100",
						 "101001010001101011101000",
						 "101001010001101010000010",
						 "101001010001101000011100",
						 "101001010001100110110110",
						 "101001010001100101010000",
						 "101001010001100011101010",
						 "101001010001100010000100",
						 "101001010001100000011110",
						 "101001010001011110111000",
						 "101001010001011101010010",
						 "101001010001011011101100",
						 "101001010001011010000110",
						 "101001010001011000100000",
						 "101001010001010110111010",
						 "101001010001010101010100",
						 "101001010001010011101110",
						 "101001010001101011110111",
						 "101001010001101010010000",
						 "101001010001101000101001",
						 "101001010001100111000010",
						 "101001010001100101011011",
						 "101001010001100011110100",
						 "101001010001100010001101",
						 "101001010001100000100110",
						 "101001010001011110111111",
						 "101001010001011101011000",
						 "101001010001011011110001",
						 "101001010001011010001010",
						 "101001010001011000100011",
						 "101001010001010110111100",
						 "101001010001010101010101",
						 "101001010001010011101110",
						 "101001010001101011110111",
						 "101001010001101010010000",
						 "101001010001101000101001",
						 "101001010001100111000010",
						 "101001010001100101011011",
						 "101001010001100011110100",
						 "101001010001100010001101",
						 "101001010001100000100110",
						 "101001010001011110111111",
						 "101001010001011101011000",
						 "101001010001011011110001",
						 "101001010001011010001010",
						 "101001010001011000100011",
						 "101001010001010110111100",
						 "101001010001010101010101",
						 "101001010001010011101110",
						 "101001010001101100000110",
						 "101001010001101010011110",
						 "101001010001101000110110",
						 "101001010001100111001110",
						 "101001010001100101100110",
						 "101001010001100011111110",
						 "101001010001100010010110",
						 "101001010001100000101110",
						 "101001010001011111000110",
						 "101001010001011101011110",
						 "101001010001011011110110",
						 "101001010001011010001110",
						 "101001010001011000100110",
						 "101001010001010110111110",
						 "101001010001010101010110",
						 "101001010001010011101110",
						 "101001010001101100000110",
						 "101001010001101010011110",
						 "101001010001101000110110",
						 "101001010001100111001110",
						 "101001010001100101100110",
						 "101001010001100011111110",
						 "101001010001100010010110",
						 "101001010001100000101110",
						 "101001010001011111000110",
						 "101001010001011101011110",
						 "101001010001011011110110",
						 "101001010001011010001110",
						 "101001010001011000100110",
						 "101001010001010110111110",
						 "101001010001010101010110",
						 "101001010001010011101110",
						 "101001010001101100000110",
						 "101001010001101010011110",
						 "101001010001101000110110",
						 "101001010001100111001110",
						 "101001010001100101100110",
						 "101001010001100011111110",
						 "101001010001100010010110",
						 "101001010001100000101110",
						 "101001010001011111000110",
						 "101001010001011101011110",
						 "101001010001011011110110",
						 "101001010001011010001110",
						 "101001010001011000100110",
						 "101001010001010110111110",
						 "101001010001010101010110",
						 "101001010001010011101110",
						 "101001001111001001010111",
						 "101001001111000111101110",
						 "101001001111000110000101",
						 "101001001111000100011100",
						 "101001001111000010110011",
						 "101001001111000001001010",
						 "101001001110111111100001",
						 "101001001110111101111000",
						 "101001001110111100001111",
						 "101001001110111010100110",
						 "101001001110111000111101",
						 "101001001110110111010100",
						 "101001001110110101101011",
						 "101001001110110100000010",
						 "101001001110110010011001",
						 "101001001110110000110000",
						 "101001001111001001010111",
						 "101001001111000111101110",
						 "101001001111000110000101",
						 "101001001111000100011100",
						 "101001001111000010110011",
						 "101001001111000001001010",
						 "101001001110111111100001",
						 "101001001110111101111000",
						 "101001001110111100001111",
						 "101001001110111010100110",
						 "101001001110111000111101",
						 "101001001110110111010100",
						 "101001001110110101101011",
						 "101001001110110100000010",
						 "101001001110110010011001",
						 "101001001110110000110000",
						 "101001001111001001010111",
						 "101001001111000111101110",
						 "101001001111000110000101",
						 "101001001111000100011100",
						 "101001001111000010110011",
						 "101001001111000001001010",
						 "101001001110111111100001",
						 "101001001110111101111000",
						 "101001001110111100001111",
						 "101001001110111010100110",
						 "101001001110111000111101",
						 "101001001110110111010100",
						 "101001001110110101101011",
						 "101001001110110100000010",
						 "101001001110110010011001",
						 "101001001110110000110000",
						 "101001001111001001100110",
						 "101001001111000111111100",
						 "101001001111000110010010",
						 "101001001111000100101000",
						 "101001001111000010111110",
						 "101001001111000001010100",
						 "101001001110111111101010",
						 "101001001110111110000000",
						 "101001001110111100010110",
						 "101001001110111010101100",
						 "101001001110111001000010",
						 "101001001110110111011000",
						 "101001001110110101101110",
						 "101001001110110100000100",
						 "101001001110110010011010",
						 "101001001110110000110000",
						 "101001001111001001100110",
						 "101001001111000111111100",
						 "101001001111000110010010",
						 "101001001111000100101000",
						 "101001001111000010111110",
						 "101001001111000001010100",
						 "101001001110111111101010",
						 "101001001110111110000000",
						 "101001001110111100010110",
						 "101001001110111010101100",
						 "101001001110111001000010",
						 "101001001110110111011000",
						 "101001001110110101101110",
						 "101001001110110100000100",
						 "101001001110110010011010",
						 "101001001110110000110000",
						 "101001001111001001100110",
						 "101001001111000111111100",
						 "101001001111000110010010",
						 "101001001111000100101000",
						 "101001001111000010111110",
						 "101001001111000001010100",
						 "101001001110111111101010",
						 "101001001110111110000000",
						 "101001001110111100010110",
						 "101001001110111010101100",
						 "101001001110111001000010",
						 "101001001110110111011000",
						 "101001001110110101101110",
						 "101001001110110100000100",
						 "101001001110110010011010",
						 "101001001110110000110000",
						 "101001001111001001110101",
						 "101001001111001000001010",
						 "101001001111000110011111",
						 "101001001111000100110100",
						 "101001001111000011001001",
						 "101001001111000001011110",
						 "101001001110111111110011",
						 "101001001110111110001000",
						 "101001001110111100011101",
						 "101001001110111010110010",
						 "101001001110111001000111",
						 "101001001110110111011100",
						 "101001001110110101110001",
						 "101001001110110100000110",
						 "101001001110110010011011",
						 "101001001110110000110000",
						 "101001001100100110110111",
						 "101001001100100101001100",
						 "101001001100100011100001",
						 "101001001100100001110110",
						 "101001001100100000001011",
						 "101001001100011110100000",
						 "101001001100011100110101",
						 "101001001100011011001010",
						 "101001001100011001011111",
						 "101001001100010111110100",
						 "101001001100010110001001",
						 "101001001100010100011110",
						 "101001001100010010110011",
						 "101001001100010001001000",
						 "101001001100001111011101",
						 "101001001100001101110010",
						 "101001001100100110110111",
						 "101001001100100101001100",
						 "101001001100100011100001",
						 "101001001100100001110110",
						 "101001001100100000001011",
						 "101001001100011110100000",
						 "101001001100011100110101",
						 "101001001100011011001010",
						 "101001001100011001011111",
						 "101001001100010111110100",
						 "101001001100010110001001",
						 "101001001100010100011110",
						 "101001001100010010110011",
						 "101001001100010001001000",
						 "101001001100001111011101",
						 "101001001100001101110010",
						 "101001001100100111000110",
						 "101001001100100101011010",
						 "101001001100100011101110",
						 "101001001100100010000010",
						 "101001001100100000010110",
						 "101001001100011110101010",
						 "101001001100011100111110",
						 "101001001100011011010010",
						 "101001001100011001100110",
						 "101001001100010111111010",
						 "101001001100010110001110",
						 "101001001100010100100010",
						 "101001001100010010110110",
						 "101001001100010001001010",
						 "101001001100001111011110",
						 "101001001100001101110010",
						 "101001001100100111000110",
						 "101001001100100101011010",
						 "101001001100100011101110",
						 "101001001100100010000010",
						 "101001001100100000010110",
						 "101001001100011110101010",
						 "101001001100011100111110",
						 "101001001100011011010010",
						 "101001001100011001100110",
						 "101001001100010111111010",
						 "101001001100010110001110",
						 "101001001100010100100010",
						 "101001001100010010110110",
						 "101001001100010001001010",
						 "101001001100001111011110",
						 "101001001100001101110010",
						 "101001001100100111000110",
						 "101001001100100101011010",
						 "101001001100100011101110",
						 "101001001100100010000010",
						 "101001001100100000010110",
						 "101001001100011110101010",
						 "101001001100011100111110",
						 "101001001100011011010010",
						 "101001001100011001100110",
						 "101001001100010111111010",
						 "101001001100010110001110",
						 "101001001100010100100010",
						 "101001001100010010110110",
						 "101001001100010001001010",
						 "101001001100001111011110",
						 "101001001100001101110010",
						 "101001001100100111010101",
						 "101001001100100101101000",
						 "101001001100100011111011",
						 "101001001100100010001110",
						 "101001001100100000100001",
						 "101001001100011110110100",
						 "101001001100011101000111",
						 "101001001100011011011010",
						 "101001001100011001101101",
						 "101001001100011000000000",
						 "101001001100010110010011",
						 "101001001100010100100110",
						 "101001001100010010111001",
						 "101001001100010001001100",
						 "101001001100001111011111",
						 "101001001100001101110010",
						 "101001001010000100010111",
						 "101001001010000010101010",
						 "101001001010000000111101",
						 "101001001001111111010000",
						 "101001001001111101100011",
						 "101001001001111011110110",
						 "101001001001111010001001",
						 "101001001001111000011100",
						 "101001001001110110101111",
						 "101001001001110101000010",
						 "101001001001110011010101",
						 "101001001001110001101000",
						 "101001001001101111111011",
						 "101001001001101110001110",
						 "101001001001101100100001",
						 "101001001001101010110100",
						 "101001001010000100100110",
						 "101001001010000010111000",
						 "101001001010000001001010",
						 "101001001001111111011100",
						 "101001001001111101101110",
						 "101001001001111100000000",
						 "101001001001111010010010",
						 "101001001001111000100100",
						 "101001001001110110110110",
						 "101001001001110101001000",
						 "101001001001110011011010",
						 "101001001001110001101100",
						 "101001001001101111111110",
						 "101001001001101110010000",
						 "101001001001101100100010",
						 "101001001001101010110100",
						 "101001001010000100100110",
						 "101001001010000010111000",
						 "101001001010000001001010",
						 "101001001001111111011100",
						 "101001001001111101101110",
						 "101001001001111100000000",
						 "101001001001111010010010",
						 "101001001001111000100100",
						 "101001001001110110110110",
						 "101001001001110101001000",
						 "101001001001110011011010",
						 "101001001001110001101100",
						 "101001001001101111111110",
						 "101001001001101110010000",
						 "101001001001101100100010",
						 "101001001001101010110100",
						 "101001001010000100100110",
						 "101001001010000010111000",
						 "101001001010000001001010",
						 "101001001001111111011100",
						 "101001001001111101101110",
						 "101001001001111100000000",
						 "101001001001111010010010",
						 "101001001001111000100100",
						 "101001001001110110110110",
						 "101001001001110101001000",
						 "101001001001110011011010",
						 "101001001001110001101100",
						 "101001001001101111111110",
						 "101001001001101110010000",
						 "101001001001101100100010",
						 "101001001001101010110100",
						 "101001001010000100110101",
						 "101001001010000011000110",
						 "101001001010000001010111",
						 "101001001001111111101000",
						 "101001001001111101111001",
						 "101001001001111100001010",
						 "101001001001111010011011",
						 "101001001001111000101100",
						 "101001001001110110111101",
						 "101001001001110101001110",
						 "101001001001110011011111",
						 "101001001001110001110000",
						 "101001001001110000000001",
						 "101001001001101110010010",
						 "101001001001101100100011",
						 "101001001001101010110100",
						 "101001001010000100110101",
						 "101001001010000011000110",
						 "101001001010000001010111",
						 "101001001001111111101000",
						 "101001001001111101111001",
						 "101001001001111100001010",
						 "101001001001111010011011",
						 "101001001001111000101100",
						 "101001001001110110111101",
						 "101001001001110101001110",
						 "101001001001110011011111",
						 "101001001001110001110000",
						 "101001001001110000000001",
						 "101001001001101110010010",
						 "101001001001101100100011",
						 "101001001001101010110100",
						 "101001000111100001110111",
						 "101001000111100000001000",
						 "101001000111011110011001",
						 "101001000111011100101010",
						 "101001000111011010111011",
						 "101001000111011001001100",
						 "101001000111010111011101",
						 "101001000111010101101110",
						 "101001000111010011111111",
						 "101001000111010010010000",
						 "101001000111010000100001",
						 "101001000111001110110010",
						 "101001000111001101000011",
						 "101001000111001011010100",
						 "101001000111001001100101",
						 "101001000111000111110110",
						 "101001000111100010000110",
						 "101001000111100000010110",
						 "101001000111011110100110",
						 "101001000111011100110110",
						 "101001000111011011000110",
						 "101001000111011001010110",
						 "101001000111010111100110",
						 "101001000111010101110110",
						 "101001000111010100000110",
						 "101001000111010010010110",
						 "101001000111010000100110",
						 "101001000111001110110110",
						 "101001000111001101000110",
						 "101001000111001011010110",
						 "101001000111001001100110",
						 "101001000111000111110110",
						 "101001000111100010000110",
						 "101001000111100000010110",
						 "101001000111011110100110",
						 "101001000111011100110110",
						 "101001000111011011000110",
						 "101001000111011001010110",
						 "101001000111010111100110",
						 "101001000111010101110110",
						 "101001000111010100000110",
						 "101001000111010010010110",
						 "101001000111010000100110",
						 "101001000111001110110110",
						 "101001000111001101000110",
						 "101001000111001011010110",
						 "101001000111001001100110",
						 "101001000111000111110110",
						 "101001000111100010000110",
						 "101001000111100000010110",
						 "101001000111011110100110",
						 "101001000111011100110110",
						 "101001000111011011000110",
						 "101001000111011001010110",
						 "101001000111010111100110",
						 "101001000111010101110110",
						 "101001000111010100000110",
						 "101001000111010010010110",
						 "101001000111010000100110",
						 "101001000111001110110110",
						 "101001000111001101000110",
						 "101001000111001011010110",
						 "101001000111001001100110",
						 "101001000111000111110110",
						 "101001000111100010010101",
						 "101001000111100000100100",
						 "101001000111011110110011",
						 "101001000111011101000010",
						 "101001000111011011010001",
						 "101001000111011001100000",
						 "101001000111010111101111",
						 "101001000111010101111110",
						 "101001000111010100001101",
						 "101001000111010010011100",
						 "101001000111010000101011",
						 "101001000111001110111010",
						 "101001000111001101001001",
						 "101001000111001011011000",
						 "101001000111001001100111",
						 "101001000111000111110110",
						 "101001000100111111010111",
						 "101001000100111101100110",
						 "101001000100111011110101",
						 "101001000100111010000100",
						 "101001000100111000010011",
						 "101001000100110110100010",
						 "101001000100110100110001",
						 "101001000100110011000000",
						 "101001000100110001001111",
						 "101001000100101111011110",
						 "101001000100101101101101",
						 "101001000100101011111100",
						 "101001000100101010001011",
						 "101001000100101000011010",
						 "101001000100100110101001",
						 "101001000100100100111000",
						 "101001000100111111010111",
						 "101001000100111101100110",
						 "101001000100111011110101",
						 "101001000100111010000100",
						 "101001000100111000010011",
						 "101001000100110110100010",
						 "101001000100110100110001",
						 "101001000100110011000000",
						 "101001000100110001001111",
						 "101001000100101111011110",
						 "101001000100101101101101",
						 "101001000100101011111100",
						 "101001000100101010001011",
						 "101001000100101000011010",
						 "101001000100100110101001",
						 "101001000100100100111000",
						 "101001000100111111100110",
						 "101001000100111101110100",
						 "101001000100111100000010",
						 "101001000100111010010000",
						 "101001000100111000011110",
						 "101001000100110110101100",
						 "101001000100110100111010",
						 "101001000100110011001000",
						 "101001000100110001010110",
						 "101001000100101111100100",
						 "101001000100101101110010",
						 "101001000100101100000000",
						 "101001000100101010001110",
						 "101001000100101000011100",
						 "101001000100100110101010",
						 "101001000100100100111000",
						 "101001000100111111100110",
						 "101001000100111101110100",
						 "101001000100111100000010",
						 "101001000100111010010000",
						 "101001000100111000011110",
						 "101001000100110110101100",
						 "101001000100110100111010",
						 "101001000100110011001000",
						 "101001000100110001010110",
						 "101001000100101111100100",
						 "101001000100101101110010",
						 "101001000100101100000000",
						 "101001000100101010001110",
						 "101001000100101000011100",
						 "101001000100100110101010",
						 "101001000100100100111000",
						 "101001000100111111100110",
						 "101001000100111101110100",
						 "101001000100111100000010",
						 "101001000100111010010000",
						 "101001000100111000011110",
						 "101001000100110110101100",
						 "101001000100110100111010",
						 "101001000100110011001000",
						 "101001000100110001010110",
						 "101001000100101111100100",
						 "101001000100101101110010",
						 "101001000100101100000000",
						 "101001000100101010001110",
						 "101001000100101000011100",
						 "101001000100100110101010",
						 "101001000100100100111000",
						 "101001000100111111110101",
						 "101001000100111110000010",
						 "101001000100111100001111",
						 "101001000100111010011100",
						 "101001000100111000101001",
						 "101001000100110110110110",
						 "101001000100110101000011",
						 "101001000100110011010000",
						 "101001000100110001011101",
						 "101001000100101111101010",
						 "101001000100101101110111",
						 "101001000100101100000100",
						 "101001000100101010010001",
						 "101001000100101000011110",
						 "101001000100100110101011",
						 "101001000100100100111000",
						 "101001000010011100110111",
						 "101001000010011011000100",
						 "101001000010011001010001",
						 "101001000010010111011110",
						 "101001000010010101101011",
						 "101001000010010011111000",
						 "101001000010010010000101",
						 "101001000010010000010010",
						 "101001000010001110011111",
						 "101001000010001100101100",
						 "101001000010001010111001",
						 "101001000010001001000110",
						 "101001000010000111010011",
						 "101001000010000101100000",
						 "101001000010000011101101",
						 "101001000010000001111010",
						 "101001000010011101000110",
						 "101001000010011011010010",
						 "101001000010011001011110",
						 "101001000010010111101010",
						 "101001000010010101110110",
						 "101001000010010100000010",
						 "101001000010010010001110",
						 "101001000010010000011010",
						 "101001000010001110100110",
						 "101001000010001100110010",
						 "101001000010001010111110",
						 "101001000010001001001010",
						 "101001000010000111010110",
						 "101001000010000101100010",
						 "101001000010000011101110",
						 "101001000010000001111010",
						 "101001000010011101000110",
						 "101001000010011011010010",
						 "101001000010011001011110",
						 "101001000010010111101010",
						 "101001000010010101110110",
						 "101001000010010100000010",
						 "101001000010010010001110",
						 "101001000010010000011010",
						 "101001000010001110100110",
						 "101001000010001100110010",
						 "101001000010001010111110",
						 "101001000010001001001010",
						 "101001000010000111010110",
						 "101001000010000101100010",
						 "101001000010000011101110",
						 "101001000010000001111010",
						 "101001000010011101000110",
						 "101001000010011011010010",
						 "101001000010011001011110",
						 "101001000010010111101010",
						 "101001000010010101110110",
						 "101001000010010100000010",
						 "101001000010010010001110",
						 "101001000010010000011010",
						 "101001000010001110100110",
						 "101001000010001100110010",
						 "101001000010001010111110",
						 "101001000010001001001010",
						 "101001000010000111010110",
						 "101001000010000101100010",
						 "101001000010000011101110",
						 "101001000010000001111010",
						 "101001000010011101010101",
						 "101001000010011011100000",
						 "101001000010011001101011",
						 "101001000010010111110110",
						 "101001000010010110000001",
						 "101001000010010100001100",
						 "101001000010010010010111",
						 "101001000010010000100010",
						 "101001000010001110101101",
						 "101001000010001100111000",
						 "101001000010001011000011",
						 "101001000010001001001110",
						 "101001000010000111011001",
						 "101001000010000101100100",
						 "101001000010000011101111",
						 "101001000010000001111010",
						 "101001000010011101010101",
						 "101001000010011011100000",
						 "101001000010011001101011",
						 "101001000010010111110110",
						 "101001000010010110000001",
						 "101001000010010100001100",
						 "101001000010010010010111",
						 "101001000010010000100010",
						 "101001000010001110101101",
						 "101001000010001100111000",
						 "101001000010001011000011",
						 "101001000010001001001110",
						 "101001000010000111011001",
						 "101001000010000101100100",
						 "101001000010000011101111",
						 "101001000010000001111010",
						 "101000111111111010010111",
						 "101000111111111000100010",
						 "101000111111110110101101",
						 "101000111111110100111000",
						 "101000111111110011000011",
						 "101000111111110001001110",
						 "101000111111101111011001",
						 "101000111111101101100100",
						 "101000111111101011101111",
						 "101000111111101001111010",
						 "101000111111101000000101",
						 "101000111111100110010000",
						 "101000111111100100011011",
						 "101000111111100010100110",
						 "101000111111100000110001",
						 "101000111111011110111100",
						 "101000111111111010100110",
						 "101000111111111000110000",
						 "101000111111110110111010",
						 "101000111111110101000100",
						 "101000111111110011001110",
						 "101000111111110001011000",
						 "101000111111101111100010",
						 "101000111111101101101100",
						 "101000111111101011110110",
						 "101000111111101010000000",
						 "101000111111101000001010",
						 "101000111111100110010100",
						 "101000111111100100011110",
						 "101000111111100010101000",
						 "101000111111100000110010",
						 "101000111111011110111100",
						 "101000111111111010100110",
						 "101000111111111000110000",
						 "101000111111110110111010",
						 "101000111111110101000100",
						 "101000111111110011001110",
						 "101000111111110001011000",
						 "101000111111101111100010",
						 "101000111111101101101100",
						 "101000111111101011110110",
						 "101000111111101010000000",
						 "101000111111101000001010",
						 "101000111111100110010100",
						 "101000111111100100011110",
						 "101000111111100010101000",
						 "101000111111100000110010",
						 "101000111111011110111100",
						 "101000111111111010100110",
						 "101000111111111000110000",
						 "101000111111110110111010",
						 "101000111111110101000100",
						 "101000111111110011001110",
						 "101000111111110001011000",
						 "101000111111101111100010",
						 "101000111111101101101100",
						 "101000111111101011110110",
						 "101000111111101010000000",
						 "101000111111101000001010",
						 "101000111111100110010100",
						 "101000111111100100011110",
						 "101000111111100010101000",
						 "101000111111100000110010",
						 "101000111111011110111100",
						 "101000111111111010110101",
						 "101000111111111000111110",
						 "101000111111110111000111",
						 "101000111111110101010000",
						 "101000111111110011011001",
						 "101000111111110001100010",
						 "101000111111101111101011",
						 "101000111111101101110100",
						 "101000111111101011111101",
						 "101000111111101010000110",
						 "101000111111101000001111",
						 "101000111111100110011000",
						 "101000111111100100100001",
						 "101000111111100010101010",
						 "101000111111100000110011",
						 "101000111111011110111100",
						 "101000111101010111110111",
						 "101000111101010110000000",
						 "101000111101010100001001",
						 "101000111101010010010010",
						 "101000111101010000011011",
						 "101000111101001110100100",
						 "101000111101001100101101",
						 "101000111101001010110110",
						 "101000111101001000111111",
						 "101000111101000111001000",
						 "101000111101000101010001",
						 "101000111101000011011010",
						 "101000111101000001100011",
						 "101000111100111111101100",
						 "101000111100111101110101",
						 "101000111100111011111110",
						 "101000111101010111110111",
						 "101000111101010110000000",
						 "101000111101010100001001",
						 "101000111101010010010010",
						 "101000111101010000011011",
						 "101000111101001110100100",
						 "101000111101001100101101",
						 "101000111101001010110110",
						 "101000111101001000111111",
						 "101000111101000111001000",
						 "101000111101000101010001",
						 "101000111101000011011010",
						 "101000111101000001100011",
						 "101000111100111111101100",
						 "101000111100111101110101",
						 "101000111100111011111110",
						 "101000111101011000000110",
						 "101000111101010110001110",
						 "101000111101010100010110",
						 "101000111101010010011110",
						 "101000111101010000100110",
						 "101000111101001110101110",
						 "101000111101001100110110",
						 "101000111101001010111110",
						 "101000111101001001000110",
						 "101000111101000111001110",
						 "101000111101000101010110",
						 "101000111101000011011110",
						 "101000111101000001100110",
						 "101000111100111111101110",
						 "101000111100111101110110",
						 "101000111100111011111110",
						 "101000111101011000000110",
						 "101000111101010110001110",
						 "101000111101010100010110",
						 "101000111101010010011110",
						 "101000111101010000100110",
						 "101000111101001110101110",
						 "101000111101001100110110",
						 "101000111101001010111110",
						 "101000111101001001000110",
						 "101000111101000111001110",
						 "101000111101000101010110",
						 "101000111101000011011110",
						 "101000111101000001100110",
						 "101000111100111111101110",
						 "101000111100111101110110",
						 "101000111100111011111110",
						 "101000111101011000000110",
						 "101000111101010110001110",
						 "101000111101010100010110",
						 "101000111101010010011110",
						 "101000111101010000100110",
						 "101000111101001110101110",
						 "101000111101001100110110",
						 "101000111101001010111110",
						 "101000111101001001000110",
						 "101000111101000111001110",
						 "101000111101000101010110",
						 "101000111101000011011110",
						 "101000111101000001100110",
						 "101000111100111111101110",
						 "101000111100111101110110",
						 "101000111100111011111110",
						 "101000111101011000010101",
						 "101000111101010110011100",
						 "101000111101010100100011",
						 "101000111101010010101010",
						 "101000111101010000110001",
						 "101000111101001110111000",
						 "101000111101001100111111",
						 "101000111101001011000110",
						 "101000111101001001001101",
						 "101000111101000111010100",
						 "101000111101000101011011",
						 "101000111101000011100010",
						 "101000111101000001101001",
						 "101000111100111111110000",
						 "101000111100111101110111",
						 "101000111100111011111110",
						 "101000111010110101010111",
						 "101000111010110011011110",
						 "101000111010110001100101",
						 "101000111010101111101100",
						 "101000111010101101110011",
						 "101000111010101011111010",
						 "101000111010101010000001",
						 "101000111010101000001000",
						 "101000111010100110001111",
						 "101000111010100100010110",
						 "101000111010100010011101",
						 "101000111010100000100100",
						 "101000111010011110101011",
						 "101000111010011100110010",
						 "101000111010011010111001",
						 "101000111010011001000000",
						 "101000111010110101010111",
						 "101000111010110011011110",
						 "101000111010110001100101",
						 "101000111010101111101100",
						 "101000111010101101110011",
						 "101000111010101011111010",
						 "101000111010101010000001",
						 "101000111010101000001000",
						 "101000111010100110001111",
						 "101000111010100100010110",
						 "101000111010100010011101",
						 "101000111010100000100100",
						 "101000111010011110101011",
						 "101000111010011100110010",
						 "101000111010011010111001",
						 "101000111010011001000000",
						 "101000111010110101100110",
						 "101000111010110011101100",
						 "101000111010110001110010",
						 "101000111010101111111000",
						 "101000111010101101111110",
						 "101000111010101100000100",
						 "101000111010101010001010",
						 "101000111010101000010000",
						 "101000111010100110010110",
						 "101000111010100100011100",
						 "101000111010100010100010",
						 "101000111010100000101000",
						 "101000111010011110101110",
						 "101000111010011100110100",
						 "101000111010011010111010",
						 "101000111010011001000000",
						 "101000111010110101100110",
						 "101000111010110011101100",
						 "101000111010110001110010",
						 "101000111010101111111000",
						 "101000111010101101111110",
						 "101000111010101100000100",
						 "101000111010101010001010",
						 "101000111010101000010000",
						 "101000111010100110010110",
						 "101000111010100100011100",
						 "101000111010100010100010",
						 "101000111010100000101000",
						 "101000111010011110101110",
						 "101000111010011100110100",
						 "101000111010011010111010",
						 "101000111010011001000000",
						 "101000111010110101100110",
						 "101000111010110011101100",
						 "101000111010110001110010",
						 "101000111010101111111000",
						 "101000111010101101111110",
						 "101000111010101100000100",
						 "101000111010101010001010",
						 "101000111010101000010000",
						 "101000111010100110010110",
						 "101000111010100100011100",
						 "101000111010100010100010",
						 "101000111010100000101000",
						 "101000111010011110101110",
						 "101000111010011100110100",
						 "101000111010011010111010",
						 "101000111010011001000000",
						 "101000111000010010110111",
						 "101000111000010000111100",
						 "101000111000001111000001",
						 "101000111000001101000110",
						 "101000111000001011001011",
						 "101000111000001001010000",
						 "101000111000000111010101",
						 "101000111000000101011010",
						 "101000111000000011011111",
						 "101000111000000001100100",
						 "101000110111111111101001",
						 "101000110111111101101110",
						 "101000110111111011110011",
						 "101000110111111001111000",
						 "101000110111110111111101",
						 "101000110111110110000010",
						 "101000111000010010110111",
						 "101000111000010000111100",
						 "101000111000001111000001",
						 "101000111000001101000110",
						 "101000111000001011001011",
						 "101000111000001001010000",
						 "101000111000000111010101",
						 "101000111000000101011010",
						 "101000111000000011011111",
						 "101000111000000001100100",
						 "101000110111111111101001",
						 "101000110111111101101110",
						 "101000110111111011110011",
						 "101000110111111001111000",
						 "101000110111110111111101",
						 "101000110111110110000010",
						 "101000111000010010110111",
						 "101000111000010000111100",
						 "101000111000001111000001",
						 "101000111000001101000110",
						 "101000111000001011001011",
						 "101000111000001001010000",
						 "101000111000000111010101",
						 "101000111000000101011010",
						 "101000111000000011011111",
						 "101000111000000001100100",
						 "101000110111111111101001",
						 "101000110111111101101110",
						 "101000110111111011110011",
						 "101000110111111001111000",
						 "101000110111110111111101",
						 "101000110111110110000010",
						 "101000111000010011000110",
						 "101000111000010001001010",
						 "101000111000001111001110",
						 "101000111000001101010010",
						 "101000111000001011010110",
						 "101000111000001001011010",
						 "101000111000000111011110",
						 "101000111000000101100010",
						 "101000111000000011100110",
						 "101000111000000001101010",
						 "101000110111111111101110",
						 "101000110111111101110010",
						 "101000110111111011110110",
						 "101000110111111001111010",
						 "101000110111110111111110",
						 "101000110111110110000010",
						 "101000111000010011000110",
						 "101000111000010001001010",
						 "101000111000001111001110",
						 "101000111000001101010010",
						 "101000111000001011010110",
						 "101000111000001001011010",
						 "101000111000000111011110",
						 "101000111000000101100010",
						 "101000111000000011100110",
						 "101000111000000001101010",
						 "101000110111111111101110",
						 "101000110111111101110010",
						 "101000110111111011110110",
						 "101000110111111001111010",
						 "101000110111110111111110",
						 "101000110111110110000010",
						 "101000110101110000001000",
						 "101000110101101110001100",
						 "101000110101101100010000",
						 "101000110101101010010100",
						 "101000110101101000011000",
						 "101000110101100110011100",
						 "101000110101100100100000",
						 "101000110101100010100100",
						 "101000110101100000101000",
						 "101000110101011110101100",
						 "101000110101011100110000",
						 "101000110101011010110100",
						 "101000110101011000111000",
						 "101000110101010110111100",
						 "101000110101010101000000",
						 "101000110101010011000100",
						 "101000110101110000010111",
						 "101000110101101110011010",
						 "101000110101101100011101",
						 "101000110101101010100000",
						 "101000110101101000100011",
						 "101000110101100110100110",
						 "101000110101100100101001",
						 "101000110101100010101100",
						 "101000110101100000101111",
						 "101000110101011110110010",
						 "101000110101011100110101",
						 "101000110101011010111000",
						 "101000110101011000111011",
						 "101000110101010110111110",
						 "101000110101010101000001",
						 "101000110101010011000100",
						 "101000110101110000010111",
						 "101000110101101110011010",
						 "101000110101101100011101",
						 "101000110101101010100000",
						 "101000110101101000100011",
						 "101000110101100110100110",
						 "101000110101100100101001",
						 "101000110101100010101100",
						 "101000110101100000101111",
						 "101000110101011110110010",
						 "101000110101011100110101",
						 "101000110101011010111000",
						 "101000110101011000111011",
						 "101000110101010110111110",
						 "101000110101010101000001",
						 "101000110101010011000100",
						 "101000110101110000100110",
						 "101000110101101110101000",
						 "101000110101101100101010",
						 "101000110101101010101100",
						 "101000110101101000101110",
						 "101000110101100110110000",
						 "101000110101100100110010",
						 "101000110101100010110100",
						 "101000110101100000110110",
						 "101000110101011110111000",
						 "101000110101011100111010",
						 "101000110101011010111100",
						 "101000110101011000111110",
						 "101000110101010111000000",
						 "101000110101010101000010",
						 "101000110101010011000100",
						 "101000110101110000100110",
						 "101000110101101110101000",
						 "101000110101101100101010",
						 "101000110101101010101100",
						 "101000110101101000101110",
						 "101000110101100110110000",
						 "101000110101100100110010",
						 "101000110101100010110100",
						 "101000110101100000110110",
						 "101000110101011110111000",
						 "101000110101011100111010",
						 "101000110101011010111100",
						 "101000110101011000111110",
						 "101000110101010111000000",
						 "101000110101010101000010",
						 "101000110101010011000100",
						 "101000110011001101101000",
						 "101000110011001011101010",
						 "101000110011001001101100",
						 "101000110011000111101110",
						 "101000110011000101110000",
						 "101000110011000011110010",
						 "101000110011000001110100",
						 "101000110010111111110110",
						 "101000110010111101111000",
						 "101000110010111011111010",
						 "101000110010111001111100",
						 "101000110010110111111110",
						 "101000110010110110000000",
						 "101000110010110100000010",
						 "101000110010110010000100",
						 "101000110010110000000110",
						 "101000110011001101110111",
						 "101000110011001011111000",
						 "101000110011001001111001",
						 "101000110011000111111010",
						 "101000110011000101111011",
						 "101000110011000011111100",
						 "101000110011000001111101",
						 "101000110010111111111110",
						 "101000110010111101111111",
						 "101000110010111100000000",
						 "101000110010111010000001",
						 "101000110010111000000010",
						 "101000110010110110000011",
						 "101000110010110100000100",
						 "101000110010110010000101",
						 "101000110010110000000110",
						 "101000110011001101110111",
						 "101000110011001011111000",
						 "101000110011001001111001",
						 "101000110011000111111010",
						 "101000110011000101111011",
						 "101000110011000011111100",
						 "101000110011000001111101",
						 "101000110010111111111110",
						 "101000110010111101111111",
						 "101000110010111100000000",
						 "101000110010111010000001",
						 "101000110010111000000010",
						 "101000110010110110000011",
						 "101000110010110100000100",
						 "101000110010110010000101",
						 "101000110010110000000110",
						 "101000110011001101110111",
						 "101000110011001011111000",
						 "101000110011001001111001",
						 "101000110011000111111010",
						 "101000110011000101111011",
						 "101000110011000011111100",
						 "101000110011000001111101",
						 "101000110010111111111110",
						 "101000110010111101111111",
						 "101000110010111100000000",
						 "101000110010111010000001",
						 "101000110010111000000010",
						 "101000110010110110000011",
						 "101000110010110100000100",
						 "101000110010110010000101",
						 "101000110010110000000110",
						 "101000110011001110000110",
						 "101000110011001100000110",
						 "101000110011001010000110",
						 "101000110011001000000110",
						 "101000110011000110000110",
						 "101000110011000100000110",
						 "101000110011000010000110",
						 "101000110011000000000110",
						 "101000110010111110000110",
						 "101000110010111100000110",
						 "101000110010111010000110",
						 "101000110010111000000110",
						 "101000110010110110000110",
						 "101000110010110100000110",
						 "101000110010110010000110",
						 "101000110010110000000110",
						 "101000110011001110000110",
						 "101000110011001100000110",
						 "101000110011001010000110",
						 "101000110011001000000110",
						 "101000110011000110000110",
						 "101000110011000100000110",
						 "101000110011000010000110",
						 "101000110011000000000110",
						 "101000110010111110000110",
						 "101000110010111100000110",
						 "101000110010111010000110",
						 "101000110010111000000110",
						 "101000110010110110000110",
						 "101000110010110100000110",
						 "101000110010110010000110",
						 "101000110010110000000110",
						 "101000110000101011001000",
						 "101000110000101001001000",
						 "101000110000100111001000",
						 "101000110000100101001000",
						 "101000110000100011001000",
						 "101000110000100001001000",
						 "101000110000011111001000",
						 "101000110000011101001000",
						 "101000110000011011001000",
						 "101000110000011001001000",
						 "101000110000010111001000",
						 "101000110000010101001000",
						 "101000110000010011001000",
						 "101000110000010001001000",
						 "101000110000001111001000",
						 "101000110000001101001000",
						 "101000110000101011010111",
						 "101000110000101001010110",
						 "101000110000100111010101",
						 "101000110000100101010100",
						 "101000110000100011010011",
						 "101000110000100001010010",
						 "101000110000011111010001",
						 "101000110000011101010000",
						 "101000110000011011001111",
						 "101000110000011001001110",
						 "101000110000010111001101",
						 "101000110000010101001100",
						 "101000110000010011001011",
						 "101000110000010001001010",
						 "101000110000001111001001",
						 "101000110000001101001000",
						 "101000110000101011010111",
						 "101000110000101001010110",
						 "101000110000100111010101",
						 "101000110000100101010100",
						 "101000110000100011010011",
						 "101000110000100001010010",
						 "101000110000011111010001",
						 "101000110000011101010000",
						 "101000110000011011001111",
						 "101000110000011001001110",
						 "101000110000010111001101",
						 "101000110000010101001100",
						 "101000110000010011001011",
						 "101000110000010001001010",
						 "101000110000001111001001",
						 "101000110000001101001000",
						 "101000110000101011010111",
						 "101000110000101001010110",
						 "101000110000100111010101",
						 "101000110000100101010100",
						 "101000110000100011010011",
						 "101000110000100001010010",
						 "101000110000011111010001",
						 "101000110000011101010000",
						 "101000110000011011001111",
						 "101000110000011001001110",
						 "101000110000010111001101",
						 "101000110000010101001100",
						 "101000110000010011001011",
						 "101000110000010001001010",
						 "101000110000001111001001",
						 "101000110000001101001000",
						 "101000110000101011100110",
						 "101000110000101001100100",
						 "101000110000100111100010",
						 "101000110000100101100000",
						 "101000110000100011011110",
						 "101000110000100001011100",
						 "101000110000011111011010",
						 "101000110000011101011000",
						 "101000110000011011010110",
						 "101000110000011001010100",
						 "101000110000010111010010",
						 "101000110000010101010000",
						 "101000110000010011001110",
						 "101000110000010001001100",
						 "101000110000001111001010",
						 "101000110000001101001000",
						 "101000101110001000101000",
						 "101000101110000110100110",
						 "101000101110000100100100",
						 "101000101110000010100010",
						 "101000101110000000100000",
						 "101000101101111110011110",
						 "101000101101111100011100",
						 "101000101101111010011010",
						 "101000101101111000011000",
						 "101000101101110110010110",
						 "101000101101110100010100",
						 "101000101101110010010010",
						 "101000101101110000010000",
						 "101000101101101110001110",
						 "101000101101101100001100",
						 "101000101101101010001010",
						 "101000101110001000101000",
						 "101000101110000110100110",
						 "101000101110000100100100",
						 "101000101110000010100010",
						 "101000101110000000100000",
						 "101000101101111110011110",
						 "101000101101111100011100",
						 "101000101101111010011010",
						 "101000101101111000011000",
						 "101000101101110110010110",
						 "101000101101110100010100",
						 "101000101101110010010010",
						 "101000101101110000010000",
						 "101000101101101110001110",
						 "101000101101101100001100",
						 "101000101101101010001010",
						 "101000101110001000110111",
						 "101000101110000110110100",
						 "101000101110000100110001",
						 "101000101110000010101110",
						 "101000101110000000101011",
						 "101000101101111110101000",
						 "101000101101111100100101",
						 "101000101101111010100010",
						 "101000101101111000011111",
						 "101000101101110110011100",
						 "101000101101110100011001",
						 "101000101101110010010110",
						 "101000101101110000010011",
						 "101000101101101110010000",
						 "101000101101101100001101",
						 "101000101101101010001010",
						 "101000101110001000110111",
						 "101000101110000110110100",
						 "101000101110000100110001",
						 "101000101110000010101110",
						 "101000101110000000101011",
						 "101000101101111110101000",
						 "101000101101111100100101",
						 "101000101101111010100010",
						 "101000101101111000011111",
						 "101000101101110110011100",
						 "101000101101110100011001",
						 "101000101101110010010110",
						 "101000101101110000010011",
						 "101000101101101110010000",
						 "101000101101101100001101",
						 "101000101101101010001010",
						 "101000101110001000110111",
						 "101000101110000110110100",
						 "101000101110000100110001",
						 "101000101110000010101110",
						 "101000101110000000101011",
						 "101000101101111110101000",
						 "101000101101111100100101",
						 "101000101101111010100010",
						 "101000101101111000011111",
						 "101000101101110110011100",
						 "101000101101110100011001",
						 "101000101101110010010110",
						 "101000101101110000010011",
						 "101000101101101110010000",
						 "101000101101101100001101",
						 "101000101101101010001010",
						 "101000101011100110001000",
						 "101000101011100100000100",
						 "101000101011100010000000",
						 "101000101011011111111100",
						 "101000101011011101111000",
						 "101000101011011011110100",
						 "101000101011011001110000",
						 "101000101011010111101100",
						 "101000101011010101101000",
						 "101000101011010011100100",
						 "101000101011010001100000",
						 "101000101011001111011100",
						 "101000101011001101011000",
						 "101000101011001011010100",
						 "101000101011001001010000",
						 "101000101011000111001100",
						 "101000101011100110001000",
						 "101000101011100100000100",
						 "101000101011100010000000",
						 "101000101011011111111100",
						 "101000101011011101111000",
						 "101000101011011011110100",
						 "101000101011011001110000",
						 "101000101011010111101100",
						 "101000101011010101101000",
						 "101000101011010011100100",
						 "101000101011010001100000",
						 "101000101011001111011100",
						 "101000101011001101011000",
						 "101000101011001011010100",
						 "101000101011001001010000",
						 "101000101011000111001100",
						 "101000101011100110001000",
						 "101000101011100100000100",
						 "101000101011100010000000",
						 "101000101011011111111100",
						 "101000101011011101111000",
						 "101000101011011011110100",
						 "101000101011011001110000",
						 "101000101011010111101100",
						 "101000101011010101101000",
						 "101000101011010011100100",
						 "101000101011010001100000",
						 "101000101011001111011100",
						 "101000101011001101011000",
						 "101000101011001011010100",
						 "101000101011001001010000",
						 "101000101011000111001100",
						 "101000101011100110010111",
						 "101000101011100100010010",
						 "101000101011100010001101",
						 "101000101011100000001000",
						 "101000101011011110000011",
						 "101000101011011011111110",
						 "101000101011011001111001",
						 "101000101011010111110100",
						 "101000101011010101101111",
						 "101000101011010011101010",
						 "101000101011010001100101",
						 "101000101011001111100000",
						 "101000101011001101011011",
						 "101000101011001011010110",
						 "101000101011001001010001",
						 "101000101011000111001100",
						 "101000101011100110010111",
						 "101000101011100100010010",
						 "101000101011100010001101",
						 "101000101011100000001000",
						 "101000101011011110000011",
						 "101000101011011011111110",
						 "101000101011011001111001",
						 "101000101011010111110100",
						 "101000101011010101101111",
						 "101000101011010011101010",
						 "101000101011010001100101",
						 "101000101011001111100000",
						 "101000101011001101011011",
						 "101000101011001011010110",
						 "101000101011001001010001",
						 "101000101011000111001100",
						 "101000101001000011011001",
						 "101000101001000001010100",
						 "101000101000111111001111",
						 "101000101000111101001010",
						 "101000101000111011000101",
						 "101000101000111001000000",
						 "101000101000110110111011",
						 "101000101000110100110110",
						 "101000101000110010110001",
						 "101000101000110000101100",
						 "101000101000101110100111",
						 "101000101000101100100010",
						 "101000101000101010011101",
						 "101000101000101000011000",
						 "101000101000100110010011",
						 "101000101000100100001110",
						 "101000101001000011101000",
						 "101000101001000001100010",
						 "101000101000111111011100",
						 "101000101000111101010110",
						 "101000101000111011010000",
						 "101000101000111001001010",
						 "101000101000110111000100",
						 "101000101000110100111110",
						 "101000101000110010111000",
						 "101000101000110000110010",
						 "101000101000101110101100",
						 "101000101000101100100110",
						 "101000101000101010100000",
						 "101000101000101000011010",
						 "101000101000100110010100",
						 "101000101000100100001110",
						 "101000101001000011101000",
						 "101000101001000001100010",
						 "101000101000111111011100",
						 "101000101000111101010110",
						 "101000101000111011010000",
						 "101000101000111001001010",
						 "101000101000110111000100",
						 "101000101000110100111110",
						 "101000101000110010111000",
						 "101000101000110000110010",
						 "101000101000101110101100",
						 "101000101000101100100110",
						 "101000101000101010100000",
						 "101000101000101000011010",
						 "101000101000100110010100",
						 "101000101000100100001110",
						 "101000101001000011101000",
						 "101000101001000001100010",
						 "101000101000111111011100",
						 "101000101000111101010110",
						 "101000101000111011010000",
						 "101000101000111001001010",
						 "101000101000110111000100",
						 "101000101000110100111110",
						 "101000101000110010111000",
						 "101000101000110000110010",
						 "101000101000101110101100",
						 "101000101000101100100110",
						 "101000101000101010100000",
						 "101000101000101000011010",
						 "101000101000100110010100",
						 "101000101000100100001110",
						 "101000100110100000111001",
						 "101000100110011110110010",
						 "101000100110011100101011",
						 "101000100110011010100100",
						 "101000100110011000011101",
						 "101000100110010110010110",
						 "101000100110010100001111",
						 "101000100110010010001000",
						 "101000100110010000000001",
						 "101000100110001101111010",
						 "101000100110001011110011",
						 "101000100110001001101100",
						 "101000100110000111100101",
						 "101000100110000101011110",
						 "101000100110000011010111",
						 "101000100110000001010000",
						 "101000100110100000111001",
						 "101000100110011110110010",
						 "101000100110011100101011",
						 "101000100110011010100100",
						 "101000100110011000011101",
						 "101000100110010110010110",
						 "101000100110010100001111",
						 "101000100110010010001000",
						 "101000100110010000000001",
						 "101000100110001101111010",
						 "101000100110001011110011",
						 "101000100110001001101100",
						 "101000100110000111100101",
						 "101000100110000101011110",
						 "101000100110000011010111",
						 "101000100110000001010000",
						 "101000100110100000111001",
						 "101000100110011110110010",
						 "101000100110011100101011",
						 "101000100110011010100100",
						 "101000100110011000011101",
						 "101000100110010110010110",
						 "101000100110010100001111",
						 "101000100110010010001000",
						 "101000100110010000000001",
						 "101000100110001101111010",
						 "101000100110001011110011",
						 "101000100110001001101100",
						 "101000100110000111100101",
						 "101000100110000101011110",
						 "101000100110000011010111",
						 "101000100110000001010000",
						 "101000100110100001001000",
						 "101000100110011111000000",
						 "101000100110011100111000",
						 "101000100110011010110000",
						 "101000100110011000101000",
						 "101000100110010110100000",
						 "101000100110010100011000",
						 "101000100110010010010000",
						 "101000100110010000001000",
						 "101000100110001110000000",
						 "101000100110001011111000",
						 "101000100110001001110000",
						 "101000100110000111101000",
						 "101000100110000101100000",
						 "101000100110000011011000",
						 "101000100110000001010000",
						 "101000100110100001001000",
						 "101000100110011111000000",
						 "101000100110011100111000",
						 "101000100110011010110000",
						 "101000100110011000101000",
						 "101000100110010110100000",
						 "101000100110010100011000",
						 "101000100110010010010000",
						 "101000100110010000001000",
						 "101000100110001110000000",
						 "101000100110001011111000",
						 "101000100110001001110000",
						 "101000100110000111101000",
						 "101000100110000101100000",
						 "101000100110000011011000",
						 "101000100110000001010000",
						 "101000100011111110001010",
						 "101000100011111100000010",
						 "101000100011111001111010",
						 "101000100011110111110010",
						 "101000100011110101101010",
						 "101000100011110011100010",
						 "101000100011110001011010",
						 "101000100011101111010010",
						 "101000100011101101001010",
						 "101000100011101011000010",
						 "101000100011101000111010",
						 "101000100011100110110010",
						 "101000100011100100101010",
						 "101000100011100010100010",
						 "101000100011100000011010",
						 "101000100011011110010010",
						 "101000100011111110011001",
						 "101000100011111100010000",
						 "101000100011111010000111",
						 "101000100011110111111110",
						 "101000100011110101110101",
						 "101000100011110011101100",
						 "101000100011110001100011",
						 "101000100011101111011010",
						 "101000100011101101010001",
						 "101000100011101011001000",
						 "101000100011101000111111",
						 "101000100011100110110110",
						 "101000100011100100101101",
						 "101000100011100010100100",
						 "101000100011100000011011",
						 "101000100011011110010010",
						 "101000100011111110011001",
						 "101000100011111100010000",
						 "101000100011111010000111",
						 "101000100011110111111110",
						 "101000100011110101110101",
						 "101000100011110011101100",
						 "101000100011110001100011",
						 "101000100011101111011010",
						 "101000100011101101010001",
						 "101000100011101011001000",
						 "101000100011101000111111",
						 "101000100011100110110110",
						 "101000100011100100101101",
						 "101000100011100010100100",
						 "101000100011100000011011",
						 "101000100011011110010010",
						 "101000100011111110011001",
						 "101000100011111100010000",
						 "101000100011111010000111",
						 "101000100011110111111110",
						 "101000100011110101110101",
						 "101000100011110011101100",
						 "101000100011110001100011",
						 "101000100011101111011010",
						 "101000100011101101010001",
						 "101000100011101011001000",
						 "101000100011101000111111",
						 "101000100011100110110110",
						 "101000100011100100101101",
						 "101000100011100010100100",
						 "101000100011100000011011",
						 "101000100011011110010010",
						 "101000100011111110101000",
						 "101000100011111100011110",
						 "101000100011111010010100",
						 "101000100011111000001010",
						 "101000100011110110000000",
						 "101000100011110011110110",
						 "101000100011110001101100",
						 "101000100011101111100010",
						 "101000100011101101011000",
						 "101000100011101011001110",
						 "101000100011101001000100",
						 "101000100011100110111010",
						 "101000100011100100110000",
						 "101000100011100010100110",
						 "101000100011100000011100",
						 "101000100011011110010010",
						 "101000100001011011101010",
						 "101000100001011001100000",
						 "101000100001010111010110",
						 "101000100001010101001100",
						 "101000100001010011000010",
						 "101000100001010000111000",
						 "101000100001001110101110",
						 "101000100001001100100100",
						 "101000100001001010011010",
						 "101000100001001000010000",
						 "101000100001000110000110",
						 "101000100001000011111100",
						 "101000100001000001110010",
						 "101000100000111111101000",
						 "101000100000111101011110",
						 "101000100000111011010100",
						 "101000100001011011101010",
						 "101000100001011001100000",
						 "101000100001010111010110",
						 "101000100001010101001100",
						 "101000100001010011000010",
						 "101000100001010000111000",
						 "101000100001001110101110",
						 "101000100001001100100100",
						 "101000100001001010011010",
						 "101000100001001000010000",
						 "101000100001000110000110",
						 "101000100001000011111100",
						 "101000100001000001110010",
						 "101000100000111111101000",
						 "101000100000111101011110",
						 "101000100000111011010100",
						 "101000100001011011111001",
						 "101000100001011001101110",
						 "101000100001010111100011",
						 "101000100001010101011000",
						 "101000100001010011001101",
						 "101000100001010001000010",
						 "101000100001001110110111",
						 "101000100001001100101100",
						 "101000100001001010100001",
						 "101000100001001000010110",
						 "101000100001000110001011",
						 "101000100001000100000000",
						 "101000100001000001110101",
						 "101000100000111111101010",
						 "101000100000111101011111",
						 "101000100000111011010100",
						 "101000100001011011111001",
						 "101000100001011001101110",
						 "101000100001010111100011",
						 "101000100001010101011000",
						 "101000100001010011001101",
						 "101000100001010001000010",
						 "101000100001001110110111",
						 "101000100001001100101100",
						 "101000100001001010100001",
						 "101000100001001000010110",
						 "101000100001000110001011",
						 "101000100001000100000000",
						 "101000100001000001110101",
						 "101000100000111111101010",
						 "101000100000111101011111",
						 "101000100000111011010100",
						 "101000100001011011111001",
						 "101000100001011001101110",
						 "101000100001010111100011",
						 "101000100001010101011000",
						 "101000100001010011001101",
						 "101000100001010001000010",
						 "101000100001001110110111",
						 "101000100001001100101100",
						 "101000100001001010100001",
						 "101000100001001000010110",
						 "101000100001000110001011",
						 "101000100001000100000000",
						 "101000100001000001110101",
						 "101000100000111111101010",
						 "101000100000111101011111",
						 "101000100000111011010100",
						 "101000011110111001001010",
						 "101000011110110110111110",
						 "101000011110110100110010",
						 "101000011110110010100110",
						 "101000011110110000011010",
						 "101000011110101110001110",
						 "101000011110101100000010",
						 "101000011110101001110110",
						 "101000011110100111101010",
						 "101000011110100101011110",
						 "101000011110100011010010",
						 "101000011110100001000110",
						 "101000011110011110111010",
						 "101000011110011100101110",
						 "101000011110011010100010",
						 "101000011110011000010110",
						 "101000011110111001001010",
						 "101000011110110110111110",
						 "101000011110110100110010",
						 "101000011110110010100110",
						 "101000011110110000011010",
						 "101000011110101110001110",
						 "101000011110101100000010",
						 "101000011110101001110110",
						 "101000011110100111101010",
						 "101000011110100101011110",
						 "101000011110100011010010",
						 "101000011110100001000110",
						 "101000011110011110111010",
						 "101000011110011100101110",
						 "101000011110011010100010",
						 "101000011110011000010110",
						 "101000011110111001001010",
						 "101000011110110110111110",
						 "101000011110110100110010",
						 "101000011110110010100110",
						 "101000011110110000011010",
						 "101000011110101110001110",
						 "101000011110101100000010",
						 "101000011110101001110110",
						 "101000011110100111101010",
						 "101000011110100101011110",
						 "101000011110100011010010",
						 "101000011110100001000110",
						 "101000011110011110111010",
						 "101000011110011100101110",
						 "101000011110011010100010",
						 "101000011110011000010110",
						 "101000011110111001011001",
						 "101000011110110111001100",
						 "101000011110110100111111",
						 "101000011110110010110010",
						 "101000011110110000100101",
						 "101000011110101110011000",
						 "101000011110101100001011",
						 "101000011110101001111110",
						 "101000011110100111110001",
						 "101000011110100101100100",
						 "101000011110100011010111",
						 "101000011110100001001010",
						 "101000011110011110111101",
						 "101000011110011100110000",
						 "101000011110011010100011",
						 "101000011110011000010110",
						 "101000011100010110011011",
						 "101000011100010100001110",
						 "101000011100010010000001",
						 "101000011100001111110100",
						 "101000011100001101100111",
						 "101000011100001011011010",
						 "101000011100001001001101",
						 "101000011100000111000000",
						 "101000011100000100110011",
						 "101000011100000010100110",
						 "101000011100000000011001",
						 "101000011011111110001100",
						 "101000011011111011111111",
						 "101000011011111001110010",
						 "101000011011110111100101",
						 "101000011011110101011000",
						 "101000011100010110011011",
						 "101000011100010100001110",
						 "101000011100010010000001",
						 "101000011100001111110100",
						 "101000011100001101100111",
						 "101000011100001011011010",
						 "101000011100001001001101",
						 "101000011100000111000000",
						 "101000011100000100110011",
						 "101000011100000010100110",
						 "101000011100000000011001",
						 "101000011011111110001100",
						 "101000011011111011111111",
						 "101000011011111001110010",
						 "101000011011110111100101",
						 "101000011011110101011000",
						 "101000011100010110101010",
						 "101000011100010100011100",
						 "101000011100010010001110",
						 "101000011100010000000000",
						 "101000011100001101110010",
						 "101000011100001011100100",
						 "101000011100001001010110",
						 "101000011100000111001000",
						 "101000011100000100111010",
						 "101000011100000010101100",
						 "101000011100000000011110",
						 "101000011011111110010000",
						 "101000011011111100000010",
						 "101000011011111001110100",
						 "101000011011110111100110",
						 "101000011011110101011000",
						 "101000011100010110101010",
						 "101000011100010100011100",
						 "101000011100010010001110",
						 "101000011100010000000000",
						 "101000011100001101110010",
						 "101000011100001011100100",
						 "101000011100001001010110",
						 "101000011100000111001000",
						 "101000011100000100111010",
						 "101000011100000010101100",
						 "101000011100000000011110",
						 "101000011011111110010000",
						 "101000011011111100000010",
						 "101000011011111001110100",
						 "101000011011110111100110",
						 "101000011011110101011000",
						 "101000011100010110101010",
						 "101000011100010100011100",
						 "101000011100010010001110",
						 "101000011100010000000000",
						 "101000011100001101110010",
						 "101000011100001011100100",
						 "101000011100001001010110",
						 "101000011100000111001000",
						 "101000011100000100111010",
						 "101000011100000010101100",
						 "101000011100000000011110",
						 "101000011011111110010000",
						 "101000011011111100000010",
						 "101000011011111001110100",
						 "101000011011110111100110",
						 "101000011011110101011000",
						 "101000011001110011101100",
						 "101000011001110001011110",
						 "101000011001101111010000",
						 "101000011001101101000010",
						 "101000011001101010110100",
						 "101000011001101000100110",
						 "101000011001100110011000",
						 "101000011001100100001010",
						 "101000011001100001111100",
						 "101000011001011111101110",
						 "101000011001011101100000",
						 "101000011001011011010010",
						 "101000011001011001000100",
						 "101000011001010110110110",
						 "101000011001010100101000",
						 "101000011001010010011010",
						 "101000011001110011111011",
						 "101000011001110001101100",
						 "101000011001101111011101",
						 "101000011001101101001110",
						 "101000011001101010111111",
						 "101000011001101000110000",
						 "101000011001100110100001",
						 "101000011001100100010010",
						 "101000011001100010000011",
						 "101000011001011111110100",
						 "101000011001011101100101",
						 "101000011001011011010110",
						 "101000011001011001000111",
						 "101000011001010110111000",
						 "101000011001010100101001",
						 "101000011001010010011010",
						 "101000011001110011111011",
						 "101000011001110001101100",
						 "101000011001101111011101",
						 "101000011001101101001110",
						 "101000011001101010111111",
						 "101000011001101000110000",
						 "101000011001100110100001",
						 "101000011001100100010010",
						 "101000011001100010000011",
						 "101000011001011111110100",
						 "101000011001011101100101",
						 "101000011001011011010110",
						 "101000011001011001000111",
						 "101000011001010110111000",
						 "101000011001010100101001",
						 "101000011001010010011010",
						 "101000011001110011111011",
						 "101000011001110001101100",
						 "101000011001101111011101",
						 "101000011001101101001110",
						 "101000011001101010111111",
						 "101000011001101000110000",
						 "101000011001100110100001",
						 "101000011001100100010010",
						 "101000011001100010000011",
						 "101000011001011111110100",
						 "101000011001011101100101",
						 "101000011001011011010110",
						 "101000011001011001000111",
						 "101000011001010110111000",
						 "101000011001010100101001",
						 "101000011001010010011010",
						 "101000010111010001001100",
						 "101000010111001110111100",
						 "101000010111001100101100",
						 "101000010111001010011100",
						 "101000010111001000001100",
						 "101000010111000101111100",
						 "101000010111000011101100",
						 "101000010111000001011100",
						 "101000010110111111001100",
						 "101000010110111100111100",
						 "101000010110111010101100",
						 "101000010110111000011100",
						 "101000010110110110001100",
						 "101000010110110011111100",
						 "101000010110110001101100",
						 "101000010110101111011100",
						 "101000010111010001001100",
						 "101000010111001110111100",
						 "101000010111001100101100",
						 "101000010111001010011100",
						 "101000010111001000001100",
						 "101000010111000101111100",
						 "101000010111000011101100",
						 "101000010111000001011100",
						 "101000010110111111001100",
						 "101000010110111100111100",
						 "101000010110111010101100",
						 "101000010110111000011100",
						 "101000010110110110001100",
						 "101000010110110011111100",
						 "101000010110110001101100",
						 "101000010110101111011100",
						 "101000010111010001001100",
						 "101000010111001110111100",
						 "101000010111001100101100",
						 "101000010111001010011100",
						 "101000010111001000001100",
						 "101000010111000101111100",
						 "101000010111000011101100",
						 "101000010111000001011100",
						 "101000010110111111001100",
						 "101000010110111100111100",
						 "101000010110111010101100",
						 "101000010110111000011100",
						 "101000010110110110001100",
						 "101000010110110011111100",
						 "101000010110110001101100",
						 "101000010110101111011100",
						 "101000010111010001011011",
						 "101000010111001111001010",
						 "101000010111001100111001",
						 "101000010111001010101000",
						 "101000010111001000010111",
						 "101000010111000110000110",
						 "101000010111000011110101",
						 "101000010111000001100100",
						 "101000010110111111010011",
						 "101000010110111101000010",
						 "101000010110111010110001",
						 "101000010110111000100000",
						 "101000010110110110001111",
						 "101000010110110011111110",
						 "101000010110110001101101",
						 "101000010110101111011100",
						 "101000010111010001011011",
						 "101000010111001111001010",
						 "101000010111001100111001",
						 "101000010111001010101000",
						 "101000010111001000010111",
						 "101000010111000110000110",
						 "101000010111000011110101",
						 "101000010111000001100100",
						 "101000010110111111010011",
						 "101000010110111101000010",
						 "101000010110111010110001",
						 "101000010110111000100000",
						 "101000010110110110001111",
						 "101000010110110011111110",
						 "101000010110110001101101",
						 "101000010110101111011100",
						 "101000010100101110011101",
						 "101000010100101100001100",
						 "101000010100101001111011",
						 "101000010100100111101010",
						 "101000010100100101011001",
						 "101000010100100011001000",
						 "101000010100100000110111",
						 "101000010100011110100110",
						 "101000010100011100010101",
						 "101000010100011010000100",
						 "101000010100010111110011",
						 "101000010100010101100010",
						 "101000010100010011010001",
						 "101000010100010001000000",
						 "101000010100001110101111",
						 "101000010100001100011110",
						 "101000010100101110101100",
						 "101000010100101100011010",
						 "101000010100101010001000",
						 "101000010100100111110110",
						 "101000010100100101100100",
						 "101000010100100011010010",
						 "101000010100100001000000",
						 "101000010100011110101110",
						 "101000010100011100011100",
						 "101000010100011010001010",
						 "101000010100010111111000",
						 "101000010100010101100110",
						 "101000010100010011010100",
						 "101000010100010001000010",
						 "101000010100001110110000",
						 "101000010100001100011110",
						 "101000010100101110101100",
						 "101000010100101100011010",
						 "101000010100101010001000",
						 "101000010100100111110110",
						 "101000010100100101100100",
						 "101000010100100011010010",
						 "101000010100100001000000",
						 "101000010100011110101110",
						 "101000010100011100011100",
						 "101000010100011010001010",
						 "101000010100010111111000",
						 "101000010100010101100110",
						 "101000010100010011010100",
						 "101000010100010001000010",
						 "101000010100001110110000",
						 "101000010100001100011110",
						 "101000010100101110101100",
						 "101000010100101100011010",
						 "101000010100101010001000",
						 "101000010100100111110110",
						 "101000010100100101100100",
						 "101000010100100011010010",
						 "101000010100100001000000",
						 "101000010100011110101110",
						 "101000010100011100011100",
						 "101000010100011010001010",
						 "101000010100010111111000",
						 "101000010100010101100110",
						 "101000010100010011010100",
						 "101000010100010001000010",
						 "101000010100001110110000",
						 "101000010100001100011110",
						 "101000010010001011111101",
						 "101000010010001001101010",
						 "101000010010000111010111",
						 "101000010010000101000100",
						 "101000010010000010110001",
						 "101000010010000000011110",
						 "101000010001111110001011",
						 "101000010001111011111000",
						 "101000010001111001100101",
						 "101000010001110111010010",
						 "101000010001110100111111",
						 "101000010001110010101100",
						 "101000010001110000011001",
						 "101000010001101110000110",
						 "101000010001101011110011",
						 "101000010001101001100000",
						 "101000010010001011111101",
						 "101000010010001001101010",
						 "101000010010000111010111",
						 "101000010010000101000100",
						 "101000010010000010110001",
						 "101000010010000000011110",
						 "101000010001111110001011",
						 "101000010001111011111000",
						 "101000010001111001100101",
						 "101000010001110111010010",
						 "101000010001110100111111",
						 "101000010001110010101100",
						 "101000010001110000011001",
						 "101000010001101110000110",
						 "101000010001101011110011",
						 "101000010001101001100000",
						 "101000010010001011111101",
						 "101000010010001001101010",
						 "101000010010000111010111",
						 "101000010010000101000100",
						 "101000010010000010110001",
						 "101000010010000000011110",
						 "101000010001111110001011",
						 "101000010001111011111000",
						 "101000010001111001100101",
						 "101000010001110111010010",
						 "101000010001110100111111",
						 "101000010001110010101100",
						 "101000010001110000011001",
						 "101000010001101110000110",
						 "101000010001101011110011",
						 "101000010001101001100000",
						 "101000010010001100001100",
						 "101000010010001001111000",
						 "101000010010000111100100",
						 "101000010010000101010000",
						 "101000010010000010111100",
						 "101000010010000000101000",
						 "101000010001111110010100",
						 "101000010001111100000000",
						 "101000010001111001101100",
						 "101000010001110111011000",
						 "101000010001110101000100",
						 "101000010001110010110000",
						 "101000010001110000011100",
						 "101000010001101110001000",
						 "101000010001101011110100",
						 "101000010001101001100000",
						 "101000010010001100001100",
						 "101000010010001001111000",
						 "101000010010000111100100",
						 "101000010010000101010000",
						 "101000010010000010111100",
						 "101000010010000000101000",
						 "101000010001111110010100",
						 "101000010001111100000000",
						 "101000010001111001101100",
						 "101000010001110111011000",
						 "101000010001110101000100",
						 "101000010001110010110000",
						 "101000010001110000011100",
						 "101000010001101110001000",
						 "101000010001101011110100",
						 "101000010001101001100000",
						 "101000001111101001001110",
						 "101000001111100110111010",
						 "101000001111100100100110",
						 "101000001111100010010010",
						 "101000001111011111111110",
						 "101000001111011101101010",
						 "101000001111011011010110",
						 "101000001111011001000010",
						 "101000001111010110101110",
						 "101000001111010100011010",
						 "101000001111010010000110",
						 "101000001111001111110010",
						 "101000001111001101011110",
						 "101000001111001011001010",
						 "101000001111001000110110",
						 "101000001111000110100010",
						 "101000001111101001011101",
						 "101000001111100111001000",
						 "101000001111100100110011",
						 "101000001111100010011110",
						 "101000001111100000001001",
						 "101000001111011101110100",
						 "101000001111011011011111",
						 "101000001111011001001010",
						 "101000001111010110110101",
						 "101000001111010100100000",
						 "101000001111010010001011",
						 "101000001111001111110110",
						 "101000001111001101100001",
						 "101000001111001011001100",
						 "101000001111001000110111",
						 "101000001111000110100010",
						 "101000001111101001011101",
						 "101000001111100111001000",
						 "101000001111100100110011",
						 "101000001111100010011110",
						 "101000001111100000001001",
						 "101000001111011101110100",
						 "101000001111011011011111",
						 "101000001111011001001010",
						 "101000001111010110110101",
						 "101000001111010100100000",
						 "101000001111010010001011",
						 "101000001111001111110110",
						 "101000001111001101100001",
						 "101000001111001011001100",
						 "101000001111001000110111",
						 "101000001111000110100010",
						 "101000001111101001011101",
						 "101000001111100111001000",
						 "101000001111100100110011",
						 "101000001111100010011110",
						 "101000001111100000001001",
						 "101000001111011101110100",
						 "101000001111011011011111",
						 "101000001111011001001010",
						 "101000001111010110110101",
						 "101000001111010100100000",
						 "101000001111010010001011",
						 "101000001111001111110110",
						 "101000001111001101100001",
						 "101000001111001011001100",
						 "101000001111001000110111",
						 "101000001111000110100010",
						 "101000001101000110101110",
						 "101000001101000100011000",
						 "101000001101000010000010",
						 "101000001100111111101100",
						 "101000001100111101010110",
						 "101000001100111011000000",
						 "101000001100111000101010",
						 "101000001100110110010100",
						 "101000001100110011111110",
						 "101000001100110001101000",
						 "101000001100101111010010",
						 "101000001100101100111100",
						 "101000001100101010100110",
						 "101000001100101000010000",
						 "101000001100100101111010",
						 "101000001100100011100100",
						 "101000001101000110101110",
						 "101000001101000100011000",
						 "101000001101000010000010",
						 "101000001100111111101100",
						 "101000001100111101010110",
						 "101000001100111011000000",
						 "101000001100111000101010",
						 "101000001100110110010100",
						 "101000001100110011111110",
						 "101000001100110001101000",
						 "101000001100101111010010",
						 "101000001100101100111100",
						 "101000001100101010100110",
						 "101000001100101000010000",
						 "101000001100100101111010",
						 "101000001100100011100100",
						 "101000001101000110101110",
						 "101000001101000100011000",
						 "101000001101000010000010",
						 "101000001100111111101100",
						 "101000001100111101010110",
						 "101000001100111011000000",
						 "101000001100111000101010",
						 "101000001100110110010100",
						 "101000001100110011111110",
						 "101000001100110001101000",
						 "101000001100101111010010",
						 "101000001100101100111100",
						 "101000001100101010100110",
						 "101000001100101000010000",
						 "101000001100100101111010",
						 "101000001100100011100100",
						 "101000001101000110101110",
						 "101000001101000100011000",
						 "101000001101000010000010",
						 "101000001100111111101100",
						 "101000001100111101010110",
						 "101000001100111011000000",
						 "101000001100111000101010",
						 "101000001100110110010100",
						 "101000001100110011111110",
						 "101000001100110001101000",
						 "101000001100101111010010",
						 "101000001100101100111100",
						 "101000001100101010100110",
						 "101000001100101000010000",
						 "101000001100100101111010",
						 "101000001100100011100100",
						 "101000001101000110111101",
						 "101000001101000100100110",
						 "101000001101000010001111",
						 "101000001100111111111000",
						 "101000001100111101100001",
						 "101000001100111011001010",
						 "101000001100111000110011",
						 "101000001100110110011100",
						 "101000001100110100000101",
						 "101000001100110001101110",
						 "101000001100101111010111",
						 "101000001100101101000000",
						 "101000001100101010101001",
						 "101000001100101000010010",
						 "101000001100100101111011",
						 "101000001100100011100100",
						 "101000001010100011111111",
						 "101000001010100001101000",
						 "101000001010011111010001",
						 "101000001010011100111010",
						 "101000001010011010100011",
						 "101000001010011000001100",
						 "101000001010010101110101",
						 "101000001010010011011110",
						 "101000001010010001000111",
						 "101000001010001110110000",
						 "101000001010001100011001",
						 "101000001010001010000010",
						 "101000001010000111101011",
						 "101000001010000101010100",
						 "101000001010000010111101",
						 "101000001010000000100110",
						 "101000001010100011111111",
						 "101000001010100001101000",
						 "101000001010011111010001",
						 "101000001010011100111010",
						 "101000001010011010100011",
						 "101000001010011000001100",
						 "101000001010010101110101",
						 "101000001010010011011110",
						 "101000001010010001000111",
						 "101000001010001110110000",
						 "101000001010001100011001",
						 "101000001010001010000010",
						 "101000001010000111101011",
						 "101000001010000101010100",
						 "101000001010000010111101",
						 "101000001010000000100110",
						 "101000001010100100001110",
						 "101000001010100001110110",
						 "101000001010011111011110",
						 "101000001010011101000110",
						 "101000001010011010101110",
						 "101000001010011000010110",
						 "101000001010010101111110",
						 "101000001010010011100110",
						 "101000001010010001001110",
						 "101000001010001110110110",
						 "101000001010001100011110",
						 "101000001010001010000110",
						 "101000001010000111101110",
						 "101000001010000101010110",
						 "101000001010000010111110",
						 "101000001010000000100110",
						 "101000001010100100001110",
						 "101000001010100001110110",
						 "101000001010011111011110",
						 "101000001010011101000110",
						 "101000001010011010101110",
						 "101000001010011000010110",
						 "101000001010010101111110",
						 "101000001010010011100110",
						 "101000001010010001001110",
						 "101000001010001110110110",
						 "101000001010001100011110",
						 "101000001010001010000110",
						 "101000001010000111101110",
						 "101000001010000101010110",
						 "101000001010000010111110",
						 "101000001010000000100110",
						 "101000001000000001010000",
						 "101000000111111110111000",
						 "101000000111111100100000",
						 "101000000111111010001000",
						 "101000000111110111110000",
						 "101000000111110101011000",
						 "101000000111110011000000",
						 "101000000111110000101000",
						 "101000000111101110010000",
						 "101000000111101011111000",
						 "101000000111101001100000",
						 "101000000111100111001000",
						 "101000000111100100110000",
						 "101000000111100010011000",
						 "101000000111100000000000",
						 "101000000111011101101000",
						 "101000001000000001011111",
						 "101000000111111111000110",
						 "101000000111111100101101",
						 "101000000111111010010100",
						 "101000000111110111111011",
						 "101000000111110101100010",
						 "101000000111110011001001",
						 "101000000111110000110000",
						 "101000000111101110010111",
						 "101000000111101011111110",
						 "101000000111101001100101",
						 "101000000111100111001100",
						 "101000000111100100110011",
						 "101000000111100010011010",
						 "101000000111100000000001",
						 "101000000111011101101000",
						 "101000001000000001011111",
						 "101000000111111111000110",
						 "101000000111111100101101",
						 "101000000111111010010100",
						 "101000000111110111111011",
						 "101000000111110101100010",
						 "101000000111110011001001",
						 "101000000111110000110000",
						 "101000000111101110010111",
						 "101000000111101011111110",
						 "101000000111101001100101",
						 "101000000111100111001100",
						 "101000000111100100110011",
						 "101000000111100010011010",
						 "101000000111100000000001",
						 "101000000111011101101000",
						 "101000001000000001011111",
						 "101000000111111111000110",
						 "101000000111111100101101",
						 "101000000111111010010100",
						 "101000000111110111111011",
						 "101000000111110101100010",
						 "101000000111110011001001",
						 "101000000111110000110000",
						 "101000000111101110010111",
						 "101000000111101011111110",
						 "101000000111101001100101",
						 "101000000111100111001100",
						 "101000000111100100110011",
						 "101000000111100010011010",
						 "101000000111100000000001",
						 "101000000111011101101000",
						 "101000000101011110110000",
						 "101000000101011100010110",
						 "101000000101011001111100",
						 "101000000101010111100010",
						 "101000000101010101001000",
						 "101000000101010010101110",
						 "101000000101010000010100",
						 "101000000101001101111010",
						 "101000000101001011100000",
						 "101000000101001001000110",
						 "101000000101000110101100",
						 "101000000101000100010010",
						 "101000000101000001111000",
						 "101000000100111111011110",
						 "101000000100111101000100",
						 "101000000100111010101010",
						 "101000000101011110110000",
						 "101000000101011100010110",
						 "101000000101011001111100",
						 "101000000101010111100010",
						 "101000000101010101001000",
						 "101000000101010010101110",
						 "101000000101010000010100",
						 "101000000101001101111010",
						 "101000000101001011100000",
						 "101000000101001001000110",
						 "101000000101000110101100",
						 "101000000101000100010010",
						 "101000000101000001111000",
						 "101000000100111111011110",
						 "101000000100111101000100",
						 "101000000100111010101010",
						 "101000000101011110110000",
						 "101000000101011100010110",
						 "101000000101011001111100",
						 "101000000101010111100010",
						 "101000000101010101001000",
						 "101000000101010010101110",
						 "101000000101010000010100",
						 "101000000101001101111010",
						 "101000000101001011100000",
						 "101000000101001001000110",
						 "101000000101000110101100",
						 "101000000101000100010010",
						 "101000000101000001111000",
						 "101000000100111111011110",
						 "101000000100111101000100",
						 "101000000100111010101010",
						 "101000000101011110111111",
						 "101000000101011100100100",
						 "101000000101011010001001",
						 "101000000101010111101110",
						 "101000000101010101010011",
						 "101000000101010010111000",
						 "101000000101010000011101",
						 "101000000101001110000010",
						 "101000000101001011100111",
						 "101000000101001001001100",
						 "101000000101000110110001",
						 "101000000101000100010110",
						 "101000000101000001111011",
						 "101000000100111111100000",
						 "101000000100111101000101",
						 "101000000100111010101010",
						 "101000000010111100000001",
						 "101000000010111001100110",
						 "101000000010110111001011",
						 "101000000010110100110000",
						 "101000000010110010010101",
						 "101000000010101111111010",
						 "101000000010101101011111",
						 "101000000010101011000100",
						 "101000000010101000101001",
						 "101000000010100110001110",
						 "101000000010100011110011",
						 "101000000010100001011000",
						 "101000000010011110111101",
						 "101000000010011100100010",
						 "101000000010011010000111",
						 "101000000010010111101100",
						 "101000000010111100000001",
						 "101000000010111001100110",
						 "101000000010110111001011",
						 "101000000010110100110000",
						 "101000000010110010010101",
						 "101000000010101111111010",
						 "101000000010101101011111",
						 "101000000010101011000100",
						 "101000000010101000101001",
						 "101000000010100110001110",
						 "101000000010100011110011",
						 "101000000010100001011000",
						 "101000000010011110111101",
						 "101000000010011100100010",
						 "101000000010011010000111",
						 "101000000010010111101100",
						 "101000000010111100000001",
						 "101000000010111001100110",
						 "101000000010110111001011",
						 "101000000010110100110000",
						 "101000000010110010010101",
						 "101000000010101111111010",
						 "101000000010101101011111",
						 "101000000010101011000100",
						 "101000000010101000101001",
						 "101000000010100110001110",
						 "101000000010100011110011",
						 "101000000010100001011000",
						 "101000000010011110111101",
						 "101000000010011100100010",
						 "101000000010011010000111",
						 "101000000010010111101100",
						 "101000000010111100010000",
						 "101000000010111001110100",
						 "101000000010110111011000",
						 "101000000010110100111100",
						 "101000000010110010100000",
						 "101000000010110000000100",
						 "101000000010101101101000",
						 "101000000010101011001100",
						 "101000000010101000110000",
						 "101000000010100110010100",
						 "101000000010100011111000",
						 "101000000010100001011100",
						 "101000000010011111000000",
						 "101000000010011100100100",
						 "101000000010011010001000",
						 "101000000010010111101100",
						 "101000000010111100010000",
						 "101000000010111001110100",
						 "101000000010110111011000",
						 "101000000010110100111100",
						 "101000000010110010100000",
						 "101000000010110000000100",
						 "101000000010101101101000",
						 "101000000010101011001100",
						 "101000000010101000110000",
						 "101000000010100110010100",
						 "101000000010100011111000",
						 "101000000010100001011100",
						 "101000000010011111000000",
						 "101000000010011100100100",
						 "101000000010011010001000",
						 "101000000010010111101100",
						 "101000000000011001010010",
						 "101000000000010110110110",
						 "101000000000010100011010",
						 "101000000000010001111110",
						 "101000000000001111100010",
						 "101000000000001101000110",
						 "101000000000001010101010",
						 "101000000000001000001110",
						 "101000000000000101110010",
						 "101000000000000011010110",
						 "101000000000000000111010",
						 "100111111111111110011110",
						 "100111111111111100000010",
						 "100111111111111001100110",
						 "100111111111110111001010",
						 "100111111111110100101110",
						 "101000000000011001100001",
						 "101000000000010111000100",
						 "101000000000010100100111",
						 "101000000000010010001010",
						 "101000000000001111101101",
						 "101000000000001101010000",
						 "101000000000001010110011",
						 "101000000000001000010110",
						 "101000000000000101111001",
						 "101000000000000011011100",
						 "101000000000000000111111",
						 "100111111111111110100010",
						 "100111111111111100000101",
						 "100111111111111001101000",
						 "100111111111110111001011",
						 "100111111111110100101110",
						 "101000000000011001100001",
						 "101000000000010111000100",
						 "101000000000010100100111",
						 "101000000000010010001010",
						 "101000000000001111101101",
						 "101000000000001101010000",
						 "101000000000001010110011",
						 "101000000000001000010110",
						 "101000000000000101111001",
						 "101000000000000011011100",
						 "101000000000000000111111",
						 "100111111111111110100010",
						 "100111111111111100000101",
						 "100111111111111001101000",
						 "100111111111110111001011",
						 "100111111111110100101110",
						 "101000000000011001100001",
						 "101000000000010111000100",
						 "101000000000010100100111",
						 "101000000000010010001010",
						 "101000000000001111101101",
						 "101000000000001101010000",
						 "101000000000001010110011",
						 "101000000000001000010110",
						 "101000000000000101111001",
						 "101000000000000011011100",
						 "101000000000000000111111",
						 "100111111111111110100010",
						 "100111111111111100000101",
						 "100111111111111001101000",
						 "100111111111110111001011",
						 "100111111111110100101110",
						 "100111111101110110110010",
						 "100111111101110100010100",
						 "100111111101110001110110",
						 "100111111101101111011000",
						 "100111111101101100111010",
						 "100111111101101010011100",
						 "100111111101100111111110",
						 "100111111101100101100000",
						 "100111111101100011000010",
						 "100111111101100000100100",
						 "100111111101011110000110",
						 "100111111101011011101000",
						 "100111111101011001001010",
						 "100111111101010110101100",
						 "100111111101010100001110",
						 "100111111101010001110000",
						 "100111111101110110110010",
						 "100111111101110100010100",
						 "100111111101110001110110",
						 "100111111101101111011000",
						 "100111111101101100111010",
						 "100111111101101010011100",
						 "100111111101100111111110",
						 "100111111101100101100000",
						 "100111111101100011000010",
						 "100111111101100000100100",
						 "100111111101011110000110",
						 "100111111101011011101000",
						 "100111111101011001001010",
						 "100111111101010110101100",
						 "100111111101010100001110",
						 "100111111101010001110000",
						 "100111111101110110110010",
						 "100111111101110100010100",
						 "100111111101110001110110",
						 "100111111101101111011000",
						 "100111111101101100111010",
						 "100111111101101010011100",
						 "100111111101100111111110",
						 "100111111101100101100000",
						 "100111111101100011000010",
						 "100111111101100000100100",
						 "100111111101011110000110",
						 "100111111101011011101000",
						 "100111111101011001001010",
						 "100111111101010110101100",
						 "100111111101010100001110",
						 "100111111101010001110000",
						 "100111111101110111000001",
						 "100111111101110100100010",
						 "100111111101110010000011",
						 "100111111101101111100100",
						 "100111111101101101000101",
						 "100111111101101010100110",
						 "100111111101101000000111",
						 "100111111101100101101000",
						 "100111111101100011001001",
						 "100111111101100000101010",
						 "100111111101011110001011",
						 "100111111101011011101100",
						 "100111111101011001001101",
						 "100111111101010110101110",
						 "100111111101010100001111",
						 "100111111101010001110000",
						 "100111111011010100000011",
						 "100111111011010001100100",
						 "100111111011001111000101",
						 "100111111011001100100110",
						 "100111111011001010000111",
						 "100111111011000111101000",
						 "100111111011000101001001",
						 "100111111011000010101010",
						 "100111111011000000001011",
						 "100111111010111101101100",
						 "100111111010111011001101",
						 "100111111010111000101110",
						 "100111111010110110001111",
						 "100111111010110011110000",
						 "100111111010110001010001",
						 "100111111010101110110010",
						 "100111111011010100000011",
						 "100111111011010001100100",
						 "100111111011001111000101",
						 "100111111011001100100110",
						 "100111111011001010000111",
						 "100111111011000111101000",
						 "100111111011000101001001",
						 "100111111011000010101010",
						 "100111111011000000001011",
						 "100111111010111101101100",
						 "100111111010111011001101",
						 "100111111010111000101110",
						 "100111111010110110001111",
						 "100111111010110011110000",
						 "100111111010110001010001",
						 "100111111010101110110010",
						 "100111111011010100000011",
						 "100111111011010001100100",
						 "100111111011001111000101",
						 "100111111011001100100110",
						 "100111111011001010000111",
						 "100111111011000111101000",
						 "100111111011000101001001",
						 "100111111011000010101010",
						 "100111111011000000001011",
						 "100111111010111101101100",
						 "100111111010111011001101",
						 "100111111010111000101110",
						 "100111111010110110001111",
						 "100111111010110011110000",
						 "100111111010110001010001",
						 "100111111010101110110010",
						 "100111111011010100010010",
						 "100111111011010001110010",
						 "100111111011001111010010",
						 "100111111011001100110010",
						 "100111111011001010010010",
						 "100111111011000111110010",
						 "100111111011000101010010",
						 "100111111011000010110010",
						 "100111111011000000010010",
						 "100111111010111101110010",
						 "100111111010111011010010",
						 "100111111010111000110010",
						 "100111111010110110010010",
						 "100111111010110011110010",
						 "100111111010110001010010",
						 "100111111010101110110010",
						 "100111111000110001010100",
						 "100111111000101110110100",
						 "100111111000101100010100",
						 "100111111000101001110100",
						 "100111111000100111010100",
						 "100111111000100100110100",
						 "100111111000100010010100",
						 "100111111000011111110100",
						 "100111111000011101010100",
						 "100111111000011010110100",
						 "100111111000011000010100",
						 "100111111000010101110100",
						 "100111111000010011010100",
						 "100111111000010000110100",
						 "100111111000001110010100",
						 "100111111000001011110100",
						 "100111111000110001010100",
						 "100111111000101110110100",
						 "100111111000101100010100",
						 "100111111000101001110100",
						 "100111111000100111010100",
						 "100111111000100100110100",
						 "100111111000100010010100",
						 "100111111000011111110100",
						 "100111111000011101010100",
						 "100111111000011010110100",
						 "100111111000011000010100",
						 "100111111000010101110100",
						 "100111111000010011010100",
						 "100111111000010000110100",
						 "100111111000001110010100",
						 "100111111000001011110100",
						 "100111111000110001100011",
						 "100111111000101111000010",
						 "100111111000101100100001",
						 "100111111000101010000000",
						 "100111111000100111011111",
						 "100111111000100100111110",
						 "100111111000100010011101",
						 "100111111000011111111100",
						 "100111111000011101011011",
						 "100111111000011010111010",
						 "100111111000011000011001",
						 "100111111000010101111000",
						 "100111111000010011010111",
						 "100111111000010000110110",
						 "100111111000001110010101",
						 "100111111000001011110100",
						 "100111111000110001100011",
						 "100111111000101111000010",
						 "100111111000101100100001",
						 "100111111000101010000000",
						 "100111111000100111011111",
						 "100111111000100100111110",
						 "100111111000100010011101",
						 "100111111000011111111100",
						 "100111111000011101011011",
						 "100111111000011010111010",
						 "100111111000011000011001",
						 "100111111000010101111000",
						 "100111111000010011010111",
						 "100111111000010000110110",
						 "100111111000001110010101",
						 "100111111000001011110100",
						 "100111110110001110100101",
						 "100111110110001100000100",
						 "100111110110001001100011",
						 "100111110110000111000010",
						 "100111110110000100100001",
						 "100111110110000010000000",
						 "100111110101111111011111",
						 "100111110101111100111110",
						 "100111110101111010011101",
						 "100111110101110111111100",
						 "100111110101110101011011",
						 "100111110101110010111010",
						 "100111110101110000011001",
						 "100111110101101101111000",
						 "100111110101101011010111",
						 "100111110101101000110110",
						 "100111110110001110110100",
						 "100111110110001100010010",
						 "100111110110001001110000",
						 "100111110110000111001110",
						 "100111110110000100101100",
						 "100111110110000010001010",
						 "100111110101111111101000",
						 "100111110101111101000110",
						 "100111110101111010100100",
						 "100111110101111000000010",
						 "100111110101110101100000",
						 "100111110101110010111110",
						 "100111110101110000011100",
						 "100111110101101101111010",
						 "100111110101101011011000",
						 "100111110101101000110110",
						 "100111110110001110110100",
						 "100111110110001100010010",
						 "100111110110001001110000",
						 "100111110110000111001110",
						 "100111110110000100101100",
						 "100111110110000010001010",
						 "100111110101111111101000",
						 "100111110101111101000110",
						 "100111110101111010100100",
						 "100111110101111000000010",
						 "100111110101110101100000",
						 "100111110101110010111110",
						 "100111110101110000011100",
						 "100111110101101101111010",
						 "100111110101101011011000",
						 "100111110101101000110110",
						 "100111110110001110110100",
						 "100111110110001100010010",
						 "100111110110001001110000",
						 "100111110110000111001110",
						 "100111110110000100101100",
						 "100111110110000010001010",
						 "100111110101111111101000",
						 "100111110101111101000110",
						 "100111110101111010100100",
						 "100111110101111000000010",
						 "100111110101110101100000",
						 "100111110101110010111110",
						 "100111110101110000011100",
						 "100111110101101101111010",
						 "100111110101101011011000",
						 "100111110101101000110110",
						 "100111110011101100000101",
						 "100111110011101001100010",
						 "100111110011100110111111",
						 "100111110011100100011100",
						 "100111110011100001111001",
						 "100111110011011111010110",
						 "100111110011011100110011",
						 "100111110011011010010000",
						 "100111110011010111101101",
						 "100111110011010101001010",
						 "100111110011010010100111",
						 "100111110011010000000100",
						 "100111110011001101100001",
						 "100111110011001010111110",
						 "100111110011001000011011",
						 "100111110011000101111000",
						 "100111110011101100000101",
						 "100111110011101001100010",
						 "100111110011100110111111",
						 "100111110011100100011100",
						 "100111110011100001111001",
						 "100111110011011111010110",
						 "100111110011011100110011",
						 "100111110011011010010000",
						 "100111110011010111101101",
						 "100111110011010101001010",
						 "100111110011010010100111",
						 "100111110011010000000100",
						 "100111110011001101100001",
						 "100111110011001010111110",
						 "100111110011001000011011",
						 "100111110011000101111000",
						 "100111110011101100000101",
						 "100111110011101001100010",
						 "100111110011100110111111",
						 "100111110011100100011100",
						 "100111110011100001111001",
						 "100111110011011111010110",
						 "100111110011011100110011",
						 "100111110011011010010000",
						 "100111110011010111101101",
						 "100111110011010101001010",
						 "100111110011010010100111",
						 "100111110011010000000100",
						 "100111110011001101100001",
						 "100111110011001010111110",
						 "100111110011001000011011",
						 "100111110011000101111000",
						 "100111110011101100000101",
						 "100111110011101001100010",
						 "100111110011100110111111",
						 "100111110011100100011100",
						 "100111110011100001111001",
						 "100111110011011111010110",
						 "100111110011011100110011",
						 "100111110011011010010000",
						 "100111110011010111101101",
						 "100111110011010101001010",
						 "100111110011010010100111",
						 "100111110011010000000100",
						 "100111110011001101100001",
						 "100111110011001010111110",
						 "100111110011001000011011",
						 "100111110011000101111000",
						 "100111110001001001010110",
						 "100111110001000110110010",
						 "100111110001000100001110",
						 "100111110001000001101010",
						 "100111110000111111000110",
						 "100111110000111100100010",
						 "100111110000111001111110",
						 "100111110000110111011010",
						 "100111110000110100110110",
						 "100111110000110010010010",
						 "100111110000101111101110",
						 "100111110000101101001010",
						 "100111110000101010100110",
						 "100111110000101000000010",
						 "100111110000100101011110",
						 "100111110000100010111010",
						 "100111110001001001010110",
						 "100111110001000110110010",
						 "100111110001000100001110",
						 "100111110001000001101010",
						 "100111110000111111000110",
						 "100111110000111100100010",
						 "100111110000111001111110",
						 "100111110000110111011010",
						 "100111110000110100110110",
						 "100111110000110010010010",
						 "100111110000101111101110",
						 "100111110000101101001010",
						 "100111110000101010100110",
						 "100111110000101000000010",
						 "100111110000100101011110",
						 "100111110000100010111010",
						 "100111110001001001010110",
						 "100111110001000110110010",
						 "100111110001000100001110",
						 "100111110001000001101010",
						 "100111110000111111000110",
						 "100111110000111100100010",
						 "100111110000111001111110",
						 "100111110000110111011010",
						 "100111110000110100110110",
						 "100111110000110010010010",
						 "100111110000101111101110",
						 "100111110000101101001010",
						 "100111110000101010100110",
						 "100111110000101000000010",
						 "100111110000100101011110",
						 "100111110000100010111010",
						 "100111110001001001100101",
						 "100111110001000111000000",
						 "100111110001000100011011",
						 "100111110001000001110110",
						 "100111110000111111010001",
						 "100111110000111100101100",
						 "100111110000111010000111",
						 "100111110000110111100010",
						 "100111110000110100111101",
						 "100111110000110010011000",
						 "100111110000101111110011",
						 "100111110000101101001110",
						 "100111110000101010101001",
						 "100111110000101000000100",
						 "100111110000100101011111",
						 "100111110000100010111010",
						 "100111101110100110100111",
						 "100111101110100100000010",
						 "100111101110100001011101",
						 "100111101110011110111000",
						 "100111101110011100010011",
						 "100111101110011001101110",
						 "100111101110010111001001",
						 "100111101110010100100100",
						 "100111101110010001111111",
						 "100111101110001111011010",
						 "100111101110001100110101",
						 "100111101110001010010000",
						 "100111101110000111101011",
						 "100111101110000101000110",
						 "100111101110000010100001",
						 "100111101101111111111100",
						 "100111101110100110100111",
						 "100111101110100100000010",
						 "100111101110100001011101",
						 "100111101110011110111000",
						 "100111101110011100010011",
						 "100111101110011001101110",
						 "100111101110010111001001",
						 "100111101110010100100100",
						 "100111101110010001111111",
						 "100111101110001111011010",
						 "100111101110001100110101",
						 "100111101110001010010000",
						 "100111101110000111101011",
						 "100111101110000101000110",
						 "100111101110000010100001",
						 "100111101101111111111100",
						 "100111101110100110110110",
						 "100111101110100100010000",
						 "100111101110100001101010",
						 "100111101110011111000100",
						 "100111101110011100011110",
						 "100111101110011001111000",
						 "100111101110010111010010",
						 "100111101110010100101100",
						 "100111101110010010000110",
						 "100111101110001111100000",
						 "100111101110001100111010",
						 "100111101110001010010100",
						 "100111101110000111101110",
						 "100111101110000101001000",
						 "100111101110000010100010",
						 "100111101101111111111100",
						 "100111101110100110110110",
						 "100111101110100100010000",
						 "100111101110100001101010",
						 "100111101110011111000100",
						 "100111101110011100011110",
						 "100111101110011001111000",
						 "100111101110010111010010",
						 "100111101110010100101100",
						 "100111101110010010000110",
						 "100111101110001111100000",
						 "100111101110001100111010",
						 "100111101110001010010100",
						 "100111101110000111101110",
						 "100111101110000101001000",
						 "100111101110000010100010",
						 "100111101101111111111100",
						 "100111101100000011111000",
						 "100111101100000001010010",
						 "100111101011111110101100",
						 "100111101011111100000110",
						 "100111101011111001100000",
						 "100111101011110110111010",
						 "100111101011110100010100",
						 "100111101011110001101110",
						 "100111101011101111001000",
						 "100111101011101100100010",
						 "100111101011101001111100",
						 "100111101011100111010110",
						 "100111101011100100110000",
						 "100111101011100010001010",
						 "100111101011011111100100",
						 "100111101011011100111110",
						 "100111101100000011111000",
						 "100111101100000001010010",
						 "100111101011111110101100",
						 "100111101011111100000110",
						 "100111101011111001100000",
						 "100111101011110110111010",
						 "100111101011110100010100",
						 "100111101011110001101110",
						 "100111101011101111001000",
						 "100111101011101100100010",
						 "100111101011101001111100",
						 "100111101011100111010110",
						 "100111101011100100110000",
						 "100111101011100010001010",
						 "100111101011011111100100",
						 "100111101011011100111110",
						 "100111101100000100000111",
						 "100111101100000001100000",
						 "100111101011111110111001",
						 "100111101011111100010010",
						 "100111101011111001101011",
						 "100111101011110111000100",
						 "100111101011110100011101",
						 "100111101011110001110110",
						 "100111101011101111001111",
						 "100111101011101100101000",
						 "100111101011101010000001",
						 "100111101011100111011010",
						 "100111101011100100110011",
						 "100111101011100010001100",
						 "100111101011011111100101",
						 "100111101011011100111110",
						 "100111101100000100000111",
						 "100111101100000001100000",
						 "100111101011111110111001",
						 "100111101011111100010010",
						 "100111101011111001101011",
						 "100111101011110111000100",
						 "100111101011110100011101",
						 "100111101011110001110110",
						 "100111101011101111001111",
						 "100111101011101100101000",
						 "100111101011101010000001",
						 "100111101011100111011010",
						 "100111101011100100110011",
						 "100111101011100010001100",
						 "100111101011011111100101",
						 "100111101011011100111110",
						 "100111101001100001001001",
						 "100111101001011110100010",
						 "100111101001011011111011",
						 "100111101001011001010100",
						 "100111101001010110101101",
						 "100111101001010100000110",
						 "100111101001010001011111",
						 "100111101001001110111000",
						 "100111101001001100010001",
						 "100111101001001001101010",
						 "100111101001000111000011",
						 "100111101001000100011100",
						 "100111101001000001110101",
						 "100111101000111111001110",
						 "100111101000111100100111",
						 "100111101000111010000000",
						 "100111101001100001011000",
						 "100111101001011110110000",
						 "100111101001011100001000",
						 "100111101001011001100000",
						 "100111101001010110111000",
						 "100111101001010100010000",
						 "100111101001010001101000",
						 "100111101001001111000000",
						 "100111101001001100011000",
						 "100111101001001001110000",
						 "100111101001000111001000",
						 "100111101001000100100000",
						 "100111101001000001111000",
						 "100111101000111111010000",
						 "100111101000111100101000",
						 "100111101000111010000000",
						 "100111101001100001011000",
						 "100111101001011110110000",
						 "100111101001011100001000",
						 "100111101001011001100000",
						 "100111101001010110111000",
						 "100111101001010100010000",
						 "100111101001010001101000",
						 "100111101001001111000000",
						 "100111101001001100011000",
						 "100111101001001001110000",
						 "100111101001000111001000",
						 "100111101001000100100000",
						 "100111101001000001111000",
						 "100111101000111111010000",
						 "100111101000111100101000",
						 "100111101000111010000000",
						 "100111101001100001011000",
						 "100111101001011110110000",
						 "100111101001011100001000",
						 "100111101001011001100000",
						 "100111101001010110111000",
						 "100111101001010100010000",
						 "100111101001010001101000",
						 "100111101001001111000000",
						 "100111101001001100011000",
						 "100111101001001001110000",
						 "100111101001000111001000",
						 "100111101001000100100000",
						 "100111101001000001111000",
						 "100111101000111111010000",
						 "100111101000111100101000",
						 "100111101000111010000000",
						 "100111100110111110011010",
						 "100111100110111011110010",
						 "100111100110111001001010",
						 "100111100110110110100010",
						 "100111100110110011111010",
						 "100111100110110001010010",
						 "100111100110101110101010",
						 "100111100110101100000010",
						 "100111100110101001011010",
						 "100111100110100110110010",
						 "100111100110100100001010",
						 "100111100110100001100010",
						 "100111100110011110111010",
						 "100111100110011100010010",
						 "100111100110011001101010",
						 "100111100110010111000010",
						 "100111100110111110101001",
						 "100111100110111100000000",
						 "100111100110111001010111",
						 "100111100110110110101110",
						 "100111100110110100000101",
						 "100111100110110001011100",
						 "100111100110101110110011",
						 "100111100110101100001010",
						 "100111100110101001100001",
						 "100111100110100110111000",
						 "100111100110100100001111",
						 "100111100110100001100110",
						 "100111100110011110111101",
						 "100111100110011100010100",
						 "100111100110011001101011",
						 "100111100110010111000010",
						 "100111100110111110101001",
						 "100111100110111100000000",
						 "100111100110111001010111",
						 "100111100110110110101110",
						 "100111100110110100000101",
						 "100111100110110001011100",
						 "100111100110101110110011",
						 "100111100110101100001010",
						 "100111100110101001100001",
						 "100111100110100110111000",
						 "100111100110100100001111",
						 "100111100110100001100110",
						 "100111100110011110111101",
						 "100111100110011100010100",
						 "100111100110011001101011",
						 "100111100110010111000010",
						 "100111100110111110101001",
						 "100111100110111100000000",
						 "100111100110111001010111",
						 "100111100110110110101110",
						 "100111100110110100000101",
						 "100111100110110001011100",
						 "100111100110101110110011",
						 "100111100110101100001010",
						 "100111100110101001100001",
						 "100111100110100110111000",
						 "100111100110100100001111",
						 "100111100110100001100110",
						 "100111100110011110111101",
						 "100111100110011100010100",
						 "100111100110011001101011",
						 "100111100110010111000010",
						 "100111100100011011111010",
						 "100111100100011001010000",
						 "100111100100010110100110",
						 "100111100100010011111100",
						 "100111100100010001010010",
						 "100111100100001110101000",
						 "100111100100001011111110",
						 "100111100100001001010100",
						 "100111100100000110101010",
						 "100111100100000100000000",
						 "100111100100000001010110",
						 "100111100011111110101100",
						 "100111100011111100000010",
						 "100111100011111001011000",
						 "100111100011110110101110",
						 "100111100011110100000100",
						 "100111100100011011111010",
						 "100111100100011001010000",
						 "100111100100010110100110",
						 "100111100100010011111100",
						 "100111100100010001010010",
						 "100111100100001110101000",
						 "100111100100001011111110",
						 "100111100100001001010100",
						 "100111100100000110101010",
						 "100111100100000100000000",
						 "100111100100000001010110",
						 "100111100011111110101100",
						 "100111100011111100000010",
						 "100111100011111001011000",
						 "100111100011110110101110",
						 "100111100011110100000100",
						 "100111100100011011111010",
						 "100111100100011001010000",
						 "100111100100010110100110",
						 "100111100100010011111100",
						 "100111100100010001010010",
						 "100111100100001110101000",
						 "100111100100001011111110",
						 "100111100100001001010100",
						 "100111100100000110101010",
						 "100111100100000100000000",
						 "100111100100000001010110",
						 "100111100011111110101100",
						 "100111100011111100000010",
						 "100111100011111001011000",
						 "100111100011110110101110",
						 "100111100011110100000100",
						 "100111100001111001001011",
						 "100111100001110110100000",
						 "100111100001110011110101",
						 "100111100001110001001010",
						 "100111100001101110011111",
						 "100111100001101011110100",
						 "100111100001101001001001",
						 "100111100001100110011110",
						 "100111100001100011110011",
						 "100111100001100001001000",
						 "100111100001011110011101",
						 "100111100001011011110010",
						 "100111100001011001000111",
						 "100111100001010110011100",
						 "100111100001010011110001",
						 "100111100001010001000110",
						 "100111100001111001001011",
						 "100111100001110110100000",
						 "100111100001110011110101",
						 "100111100001110001001010",
						 "100111100001101110011111",
						 "100111100001101011110100",
						 "100111100001101001001001",
						 "100111100001100110011110",
						 "100111100001100011110011",
						 "100111100001100001001000",
						 "100111100001011110011101",
						 "100111100001011011110010",
						 "100111100001011001000111",
						 "100111100001010110011100",
						 "100111100001010011110001",
						 "100111100001010001000110",
						 "100111100001111001001011",
						 "100111100001110110100000",
						 "100111100001110011110101",
						 "100111100001110001001010",
						 "100111100001101110011111",
						 "100111100001101011110100",
						 "100111100001101001001001",
						 "100111100001100110011110",
						 "100111100001100011110011",
						 "100111100001100001001000",
						 "100111100001011110011101",
						 "100111100001011011110010",
						 "100111100001011001000111",
						 "100111100001010110011100",
						 "100111100001010011110001",
						 "100111100001010001000110",
						 "100111100001111001001011",
						 "100111100001110110100000",
						 "100111100001110011110101",
						 "100111100001110001001010",
						 "100111100001101110011111",
						 "100111100001101011110100",
						 "100111100001101001001001",
						 "100111100001100110011110",
						 "100111100001100011110011",
						 "100111100001100001001000",
						 "100111100001011110011101",
						 "100111100001011011110010",
						 "100111100001011001000111",
						 "100111100001010110011100",
						 "100111100001010011110001",
						 "100111100001010001000110",
						 "100111011111010110011100",
						 "100111011111010011110000",
						 "100111011111010001000100",
						 "100111011111001110011000",
						 "100111011111001011101100",
						 "100111011111001001000000",
						 "100111011111000110010100",
						 "100111011111000011101000",
						 "100111011111000000111100",
						 "100111011110111110010000",
						 "100111011110111011100100",
						 "100111011110111000111000",
						 "100111011110110110001100",
						 "100111011110110011100000",
						 "100111011110110000110100",
						 "100111011110101110001000",
						 "100111011111010110011100",
						 "100111011111010011110000",
						 "100111011111010001000100",
						 "100111011111001110011000",
						 "100111011111001011101100",
						 "100111011111001001000000",
						 "100111011111000110010100",
						 "100111011111000011101000",
						 "100111011111000000111100",
						 "100111011110111110010000",
						 "100111011110111011100100",
						 "100111011110111000111000",
						 "100111011110110110001100",
						 "100111011110110011100000",
						 "100111011110110000110100",
						 "100111011110101110001000",
						 "100111011111010110011100",
						 "100111011111010011110000",
						 "100111011111010001000100",
						 "100111011111001110011000",
						 "100111011111001011101100",
						 "100111011111001001000000",
						 "100111011111000110010100",
						 "100111011111000011101000",
						 "100111011111000000111100",
						 "100111011110111110010000",
						 "100111011110111011100100",
						 "100111011110111000111000",
						 "100111011110110110001100",
						 "100111011110110011100000",
						 "100111011110110000110100",
						 "100111011110101110001000",
						 "100111011111010110101011",
						 "100111011111010011111110",
						 "100111011111010001010001",
						 "100111011111001110100100",
						 "100111011111001011110111",
						 "100111011111001001001010",
						 "100111011111000110011101",
						 "100111011111000011110000",
						 "100111011111000001000011",
						 "100111011110111110010110",
						 "100111011110111011101001",
						 "100111011110111000111100",
						 "100111011110110110001111",
						 "100111011110110011100010",
						 "100111011110110000110101",
						 "100111011110101110001000",
						 "100111011100110011101101",
						 "100111011100110001000000",
						 "100111011100101110010011",
						 "100111011100101011100110",
						 "100111011100101000111001",
						 "100111011100100110001100",
						 "100111011100100011011111",
						 "100111011100100000110010",
						 "100111011100011110000101",
						 "100111011100011011011000",
						 "100111011100011000101011",
						 "100111011100010101111110",
						 "100111011100010011010001",
						 "100111011100010000100100",
						 "100111011100001101110111",
						 "100111011100001011001010",
						 "100111011100110011101101",
						 "100111011100110001000000",
						 "100111011100101110010011",
						 "100111011100101011100110",
						 "100111011100101000111001",
						 "100111011100100110001100",
						 "100111011100100011011111",
						 "100111011100100000110010",
						 "100111011100011110000101",
						 "100111011100011011011000",
						 "100111011100011000101011",
						 "100111011100010101111110",
						 "100111011100010011010001",
						 "100111011100010000100100",
						 "100111011100001101110111",
						 "100111011100001011001010",
						 "100111011100110011101101",
						 "100111011100110001000000",
						 "100111011100101110010011",
						 "100111011100101011100110",
						 "100111011100101000111001",
						 "100111011100100110001100",
						 "100111011100100011011111",
						 "100111011100100000110010",
						 "100111011100011110000101",
						 "100111011100011011011000",
						 "100111011100011000101011",
						 "100111011100010101111110",
						 "100111011100010011010001",
						 "100111011100010000100100",
						 "100111011100001101110111",
						 "100111011100001011001010",
						 "100111011100110011111100",
						 "100111011100110001001110",
						 "100111011100101110100000",
						 "100111011100101011110010",
						 "100111011100101001000100",
						 "100111011100100110010110",
						 "100111011100100011101000",
						 "100111011100100000111010",
						 "100111011100011110001100",
						 "100111011100011011011110",
						 "100111011100011000110000",
						 "100111011100010110000010",
						 "100111011100010011010100",
						 "100111011100010000100110",
						 "100111011100001101111000",
						 "100111011100001011001010",
						 "100111011010010000111110",
						 "100111011010001110010000",
						 "100111011010001011100010",
						 "100111011010001000110100",
						 "100111011010000110000110",
						 "100111011010000011011000",
						 "100111011010000000101010",
						 "100111011001111101111100",
						 "100111011001111011001110",
						 "100111011001111000100000",
						 "100111011001110101110010",
						 "100111011001110011000100",
						 "100111011001110000010110",
						 "100111011001101101101000",
						 "100111011001101010111010",
						 "100111011001101000001100",
						 "100111011010010000111110",
						 "100111011010001110010000",
						 "100111011010001011100010",
						 "100111011010001000110100",
						 "100111011010000110000110",
						 "100111011010000011011000",
						 "100111011010000000101010",
						 "100111011001111101111100",
						 "100111011001111011001110",
						 "100111011001111000100000",
						 "100111011001110101110010",
						 "100111011001110011000100",
						 "100111011001110000010110",
						 "100111011001101101101000",
						 "100111011001101010111010",
						 "100111011001101000001100",
						 "100111011010010001001101",
						 "100111011010001110011110",
						 "100111011010001011101111",
						 "100111011010001001000000",
						 "100111011010000110010001",
						 "100111011010000011100010",
						 "100111011010000000110011",
						 "100111011001111110000100",
						 "100111011001111011010101",
						 "100111011001111000100110",
						 "100111011001110101110111",
						 "100111011001110011001000",
						 "100111011001110000011001",
						 "100111011001101101101010",
						 "100111011001101010111011",
						 "100111011001101000001100",
						 "100111010111101110001111",
						 "100111010111101011100000",
						 "100111010111101000110001",
						 "100111010111100110000010",
						 "100111010111100011010011",
						 "100111010111100000100100",
						 "100111010111011101110101",
						 "100111010111011011000110",
						 "100111010111011000010111",
						 "100111010111010101101000",
						 "100111010111010010111001",
						 "100111010111010000001010",
						 "100111010111001101011011",
						 "100111010111001010101100",
						 "100111010111000111111101",
						 "100111010111000101001110",
						 "100111010111101110001111",
						 "100111010111101011100000",
						 "100111010111101000110001",
						 "100111010111100110000010",
						 "100111010111100011010011",
						 "100111010111100000100100",
						 "100111010111011101110101",
						 "100111010111011011000110",
						 "100111010111011000010111",
						 "100111010111010101101000",
						 "100111010111010010111001",
						 "100111010111010000001010",
						 "100111010111001101011011",
						 "100111010111001010101100",
						 "100111010111000111111101",
						 "100111010111000101001110",
						 "100111010111101110001111",
						 "100111010111101011100000",
						 "100111010111101000110001",
						 "100111010111100110000010",
						 "100111010111100011010011",
						 "100111010111100000100100",
						 "100111010111011101110101",
						 "100111010111011011000110",
						 "100111010111011000010111",
						 "100111010111010101101000",
						 "100111010111010010111001",
						 "100111010111010000001010",
						 "100111010111001101011011",
						 "100111010111001010101100",
						 "100111010111000111111101",
						 "100111010111000101001110",
						 "100111010111101110011110",
						 "100111010111101011101110",
						 "100111010111101000111110",
						 "100111010111100110001110",
						 "100111010111100011011110",
						 "100111010111100000101110",
						 "100111010111011101111110",
						 "100111010111011011001110",
						 "100111010111011000011110",
						 "100111010111010101101110",
						 "100111010111010010111110",
						 "100111010111010000001110",
						 "100111010111001101011110",
						 "100111010111001010101110",
						 "100111010111000111111110",
						 "100111010111000101001110",
						 "100111010101001011100000",
						 "100111010101001000110000",
						 "100111010101000110000000",
						 "100111010101000011010000",
						 "100111010101000000100000",
						 "100111010100111101110000",
						 "100111010100111011000000",
						 "100111010100111000010000",
						 "100111010100110101100000",
						 "100111010100110010110000",
						 "100111010100110000000000",
						 "100111010100101101010000",
						 "100111010100101010100000",
						 "100111010100100111110000",
						 "100111010100100101000000",
						 "100111010100100010010000",
						 "100111010101001011100000",
						 "100111010101001000110000",
						 "100111010101000110000000",
						 "100111010101000011010000",
						 "100111010101000000100000",
						 "100111010100111101110000",
						 "100111010100111011000000",
						 "100111010100111000010000",
						 "100111010100110101100000",
						 "100111010100110010110000",
						 "100111010100110000000000",
						 "100111010100101101010000",
						 "100111010100101010100000",
						 "100111010100100111110000",
						 "100111010100100101000000",
						 "100111010100100010010000",
						 "100111010101001011101111",
						 "100111010101001000111110",
						 "100111010101000110001101",
						 "100111010101000011011100",
						 "100111010101000000101011",
						 "100111010100111101111010",
						 "100111010100111011001001",
						 "100111010100111000011000",
						 "100111010100110101100111",
						 "100111010100110010110110",
						 "100111010100110000000101",
						 "100111010100101101010100",
						 "100111010100101010100011",
						 "100111010100100111110010",
						 "100111010100100101000001",
						 "100111010100100010010000",
						 "100111010101001011101111",
						 "100111010101001000111110",
						 "100111010101000110001101",
						 "100111010101000011011100",
						 "100111010101000000101011",
						 "100111010100111101111010",
						 "100111010100111011001001",
						 "100111010100111000011000",
						 "100111010100110101100111",
						 "100111010100110010110110",
						 "100111010100110000000101",
						 "100111010100101101010100",
						 "100111010100101010100011",
						 "100111010100100111110010",
						 "100111010100100101000001",
						 "100111010100100010010000",
						 "100111010010101000110001",
						 "100111010010100110000000",
						 "100111010010100011001111",
						 "100111010010100000011110",
						 "100111010010011101101101",
						 "100111010010011010111100",
						 "100111010010011000001011",
						 "100111010010010101011010",
						 "100111010010010010101001",
						 "100111010010001111111000",
						 "100111010010001101000111",
						 "100111010010001010010110",
						 "100111010010000111100101",
						 "100111010010000100110100",
						 "100111010010000010000011",
						 "100111010001111111010010",
						 "100111010010101000110001",
						 "100111010010100110000000",
						 "100111010010100011001111",
						 "100111010010100000011110",
						 "100111010010011101101101",
						 "100111010010011010111100",
						 "100111010010011000001011",
						 "100111010010010101011010",
						 "100111010010010010101001",
						 "100111010010001111111000",
						 "100111010010001101000111",
						 "100111010010001010010110",
						 "100111010010000111100101",
						 "100111010010000100110100",
						 "100111010010000010000011",
						 "100111010001111111010010",
						 "100111010010101001000000",
						 "100111010010100110001110",
						 "100111010010100011011100",
						 "100111010010100000101010",
						 "100111010010011101111000",
						 "100111010010011011000110",
						 "100111010010011000010100",
						 "100111010010010101100010",
						 "100111010010010010110000",
						 "100111010010001111111110",
						 "100111010010001101001100",
						 "100111010010001010011010",
						 "100111010010000111101000",
						 "100111010010000100110110",
						 "100111010010000010000100",
						 "100111010001111111010010",
						 "100111010010101001000000",
						 "100111010010100110001110",
						 "100111010010100011011100",
						 "100111010010100000101010",
						 "100111010010011101111000",
						 "100111010010011011000110",
						 "100111010010011000010100",
						 "100111010010010101100010",
						 "100111010010010010110000",
						 "100111010010001111111110",
						 "100111010010001101001100",
						 "100111010010001010011010",
						 "100111010010000111101000",
						 "100111010010000100110110",
						 "100111010010000010000100",
						 "100111010001111111010010",
						 "100111010000000110000010",
						 "100111010000000011010000",
						 "100111010000000000011110",
						 "100111001111111101101100",
						 "100111001111111010111010",
						 "100111001111111000001000",
						 "100111001111110101010110",
						 "100111001111110010100100",
						 "100111001111101111110010",
						 "100111001111101101000000",
						 "100111001111101010001110",
						 "100111001111100111011100",
						 "100111001111100100101010",
						 "100111001111100001111000",
						 "100111001111011111000110",
						 "100111001111011100010100",
						 "100111010000000110010001",
						 "100111010000000011011110",
						 "100111010000000000101011",
						 "100111001111111101111000",
						 "100111001111111011000101",
						 "100111001111111000010010",
						 "100111001111110101011111",
						 "100111001111110010101100",
						 "100111001111101111111001",
						 "100111001111101101000110",
						 "100111001111101010010011",
						 "100111001111100111100000",
						 "100111001111100100101101",
						 "100111001111100001111010",
						 "100111001111011111000111",
						 "100111001111011100010100",
						 "100111010000000110010001",
						 "100111010000000011011110",
						 "100111010000000000101011",
						 "100111001111111101111000",
						 "100111001111111011000101",
						 "100111001111111000010010",
						 "100111001111110101011111",
						 "100111001111110010101100",
						 "100111001111101111111001",
						 "100111001111101101000110",
						 "100111001111101010010011",
						 "100111001111100111100000",
						 "100111001111100100101101",
						 "100111001111100001111010",
						 "100111001111011111000111",
						 "100111001111011100010100",
						 "100111001101100011010011",
						 "100111001101100000100000",
						 "100111001101011101101101",
						 "100111001101011010111010",
						 "100111001101011000000111",
						 "100111001101010101010100",
						 "100111001101010010100001",
						 "100111001101001111101110",
						 "100111001101001100111011",
						 "100111001101001010001000",
						 "100111001101000111010101",
						 "100111001101000100100010",
						 "100111001101000001101111",
						 "100111001100111110111100",
						 "100111001100111100001001",
						 "100111001100111001010110",
						 "100111001101100011010011",
						 "100111001101100000100000",
						 "100111001101011101101101",
						 "100111001101011010111010",
						 "100111001101011000000111",
						 "100111001101010101010100",
						 "100111001101010010100001",
						 "100111001101001111101110",
						 "100111001101001100111011",
						 "100111001101001010001000",
						 "100111001101000111010101",
						 "100111001101000100100010",
						 "100111001101000001101111",
						 "100111001100111110111100",
						 "100111001100111100001001",
						 "100111001100111001010110",
						 "100111001101100011100010",
						 "100111001101100000101110",
						 "100111001101011101111010",
						 "100111001101011011000110",
						 "100111001101011000010010",
						 "100111001101010101011110",
						 "100111001101010010101010",
						 "100111001101001111110110",
						 "100111001101001101000010",
						 "100111001101001010001110",
						 "100111001101000111011010",
						 "100111001101000100100110",
						 "100111001101000001110010",
						 "100111001100111110111110",
						 "100111001100111100001010",
						 "100111001100111001010110",
						 "100111001101100011100010",
						 "100111001101100000101110",
						 "100111001101011101111010",
						 "100111001101011011000110",
						 "100111001101011000010010",
						 "100111001101010101011110",
						 "100111001101010010101010",
						 "100111001101001111110110",
						 "100111001101001101000010",
						 "100111001101001010001110",
						 "100111001101000111011010",
						 "100111001101000100100110",
						 "100111001101000001110010",
						 "100111001100111110111110",
						 "100111001100111100001010",
						 "100111001100111001010110",
						 "100111001011000000100100",
						 "100111001010111101110000",
						 "100111001010111010111100",
						 "100111001010111000001000",
						 "100111001010110101010100",
						 "100111001010110010100000",
						 "100111001010101111101100",
						 "100111001010101100111000",
						 "100111001010101010000100",
						 "100111001010100111010000",
						 "100111001010100100011100",
						 "100111001010100001101000",
						 "100111001010011110110100",
						 "100111001010011100000000",
						 "100111001010011001001100",
						 "100111001010010110011000",
						 "100111001011000000100100",
						 "100111001010111101110000",
						 "100111001010111010111100",
						 "100111001010111000001000",
						 "100111001010110101010100",
						 "100111001010110010100000",
						 "100111001010101111101100",
						 "100111001010101100111000",
						 "100111001010101010000100",
						 "100111001010100111010000",
						 "100111001010100100011100",
						 "100111001010100001101000",
						 "100111001010011110110100",
						 "100111001010011100000000",
						 "100111001010011001001100",
						 "100111001010010110011000",
						 "100111001011000000110011",
						 "100111001010111101111110",
						 "100111001010111011001001",
						 "100111001010111000010100",
						 "100111001010110101011111",
						 "100111001010110010101010",
						 "100111001010101111110101",
						 "100111001010101101000000",
						 "100111001010101010001011",
						 "100111001010100111010110",
						 "100111001010100100100001",
						 "100111001010100001101100",
						 "100111001010011110110111",
						 "100111001010011100000010",
						 "100111001010011001001101",
						 "100111001010010110011000",
						 "100111001000011101110101",
						 "100111001000011011000000",
						 "100111001000011000001011",
						 "100111001000010101010110",
						 "100111001000010010100001",
						 "100111001000001111101100",
						 "100111001000001100110111",
						 "100111001000001010000010",
						 "100111001000000111001101",
						 "100111001000000100011000",
						 "100111001000000001100011",
						 "100111000111111110101110",
						 "100111000111111011111001",
						 "100111000111111001000100",
						 "100111000111110110001111",
						 "100111000111110011011010",
						 "100111001000011101110101",
						 "100111001000011011000000",
						 "100111001000011000001011",
						 "100111001000010101010110",
						 "100111001000010010100001",
						 "100111001000001111101100",
						 "100111001000001100110111",
						 "100111001000001010000010",
						 "100111001000000111001101",
						 "100111001000000100011000",
						 "100111001000000001100011",
						 "100111000111111110101110",
						 "100111000111111011111001",
						 "100111000111111001000100",
						 "100111000111110110001111",
						 "100111000111110011011010",
						 "100111001000011110000100",
						 "100111001000011011001110",
						 "100111001000011000011000",
						 "100111001000010101100010",
						 "100111001000010010101100",
						 "100111001000001111110110",
						 "100111001000001101000000",
						 "100111001000001010001010",
						 "100111001000000111010100",
						 "100111001000000100011110",
						 "100111001000000001101000",
						 "100111000111111110110010",
						 "100111000111111011111100",
						 "100111000111111001000110",
						 "100111000111110110010000",
						 "100111000111110011011010",
						 "100111001000011110000100",
						 "100111001000011011001110",
						 "100111001000011000011000",
						 "100111001000010101100010",
						 "100111001000010010101100",
						 "100111001000001111110110",
						 "100111001000001101000000",
						 "100111001000001010001010",
						 "100111001000000111010100",
						 "100111001000000100011110",
						 "100111001000000001101000",
						 "100111000111111110110010",
						 "100111000111111011111100",
						 "100111000111111001000110",
						 "100111000111110110010000",
						 "100111000111110011011010",
						 "100111000101111011000110",
						 "100111000101111000010000",
						 "100111000101110101011010",
						 "100111000101110010100100",
						 "100111000101101111101110",
						 "100111000101101100111000",
						 "100111000101101010000010",
						 "100111000101100111001100",
						 "100111000101100100010110",
						 "100111000101100001100000",
						 "100111000101011110101010",
						 "100111000101011011110100",
						 "100111000101011000111110",
						 "100111000101010110001000",
						 "100111000101010011010010",
						 "100111000101010000011100",
						 "100111000101111011000110",
						 "100111000101111000010000",
						 "100111000101110101011010",
						 "100111000101110010100100",
						 "100111000101101111101110",
						 "100111000101101100111000",
						 "100111000101101010000010",
						 "100111000101100111001100",
						 "100111000101100100010110",
						 "100111000101100001100000",
						 "100111000101011110101010",
						 "100111000101011011110100",
						 "100111000101011000111110",
						 "100111000101010110001000",
						 "100111000101010011010010",
						 "100111000101010000011100",
						 "100111000101111011010101",
						 "100111000101111000011110",
						 "100111000101110101100111",
						 "100111000101110010110000",
						 "100111000101101111111001",
						 "100111000101101101000010",
						 "100111000101101010001011",
						 "100111000101100111010100",
						 "100111000101100100011101",
						 "100111000101100001100110",
						 "100111000101011110101111",
						 "100111000101011011111000",
						 "100111000101011001000001",
						 "100111000101010110001010",
						 "100111000101010011010011",
						 "100111000101010000011100",
						 "100111000101111011010101",
						 "100111000101111000011110",
						 "100111000101110101100111",
						 "100111000101110010110000",
						 "100111000101101111111001",
						 "100111000101101101000010",
						 "100111000101101010001011",
						 "100111000101100111010100",
						 "100111000101100100011101",
						 "100111000101100001100110",
						 "100111000101011110101111",
						 "100111000101011011111000",
						 "100111000101011001000001",
						 "100111000101010110001010",
						 "100111000101010011010011",
						 "100111000101010000011100",
						 "100111000011011000010111",
						 "100111000011010101100000",
						 "100111000011010010101001",
						 "100111000011001111110010",
						 "100111000011001100111011",
						 "100111000011001010000100",
						 "100111000011000111001101",
						 "100111000011000100010110",
						 "100111000011000001011111",
						 "100111000010111110101000",
						 "100111000010111011110001",
						 "100111000010111000111010",
						 "100111000010110110000011",
						 "100111000010110011001100",
						 "100111000010110000010101",
						 "100111000010101101011110",
						 "100111000011011000010111",
						 "100111000011010101100000",
						 "100111000011010010101001",
						 "100111000011001111110010",
						 "100111000011001100111011",
						 "100111000011001010000100",
						 "100111000011000111001101",
						 "100111000011000100010110",
						 "100111000011000001011111",
						 "100111000010111110101000",
						 "100111000010111011110001",
						 "100111000010111000111010",
						 "100111000010110110000011",
						 "100111000010110011001100",
						 "100111000010110000010101",
						 "100111000010101101011110",
						 "100111000011011000100110",
						 "100111000011010101101110",
						 "100111000011010010110110",
						 "100111000011001111111110",
						 "100111000011001101000110",
						 "100111000011001010001110",
						 "100111000011000111010110",
						 "100111000011000100011110",
						 "100111000011000001100110",
						 "100111000010111110101110",
						 "100111000010111011110110",
						 "100111000010111000111110",
						 "100111000010110110000110",
						 "100111000010110011001110",
						 "100111000010110000010110",
						 "100111000010101101011110",
						 "100111000000110101101000",
						 "100111000000110010110000",
						 "100111000000101111111000",
						 "100111000000101101000000",
						 "100111000000101010001000",
						 "100111000000100111010000",
						 "100111000000100100011000",
						 "100111000000100001100000",
						 "100111000000011110101000",
						 "100111000000011011110000",
						 "100111000000011000111000",
						 "100111000000010110000000",
						 "100111000000010011001000",
						 "100111000000010000010000",
						 "100111000000001101011000",
						 "100111000000001010100000",
						 "100111000000110101101000",
						 "100111000000110010110000",
						 "100111000000101111111000",
						 "100111000000101101000000",
						 "100111000000101010001000",
						 "100111000000100111010000",
						 "100111000000100100011000",
						 "100111000000100001100000",
						 "100111000000011110101000",
						 "100111000000011011110000",
						 "100111000000011000111000",
						 "100111000000010110000000",
						 "100111000000010011001000",
						 "100111000000010000010000",
						 "100111000000001101011000",
						 "100111000000001010100000",
						 "100111000000110101110111",
						 "100111000000110010111110",
						 "100111000000110000000101",
						 "100111000000101101001100",
						 "100111000000101010010011",
						 "100111000000100111011010",
						 "100111000000100100100001",
						 "100111000000100001101000",
						 "100111000000011110101111",
						 "100111000000011011110110",
						 "100111000000011000111101",
						 "100111000000010110000100",
						 "100111000000010011001011",
						 "100111000000010000010010",
						 "100111000000001101011001",
						 "100111000000001010100000",
						 "100111000000110101110111",
						 "100111000000110010111110",
						 "100111000000110000000101",
						 "100111000000101101001100",
						 "100111000000101010010011",
						 "100111000000100111011010",
						 "100111000000100100100001",
						 "100111000000100001101000",
						 "100111000000011110101111",
						 "100111000000011011110110",
						 "100111000000011000111101",
						 "100111000000010110000100",
						 "100111000000010011001011",
						 "100111000000010000010010",
						 "100111000000001101011001",
						 "100111000000001010100000",
						 "100110111110010010111001",
						 "100110111110010000000000",
						 "100110111110001101000111",
						 "100110111110001010001110",
						 "100110111110000111010101",
						 "100110111110000100011100",
						 "100110111110000001100011",
						 "100110111101111110101010",
						 "100110111101111011110001",
						 "100110111101111000111000",
						 "100110111101110101111111",
						 "100110111101110011000110",
						 "100110111101110000001101",
						 "100110111101101101010100",
						 "100110111101101010011011",
						 "100110111101100111100010",
						 "100110111110010010111001",
						 "100110111110010000000000",
						 "100110111110001101000111",
						 "100110111110001010001110",
						 "100110111110000111010101",
						 "100110111110000100011100",
						 "100110111110000001100011",
						 "100110111101111110101010",
						 "100110111101111011110001",
						 "100110111101111000111000",
						 "100110111101110101111111",
						 "100110111101110011000110",
						 "100110111101110000001101",
						 "100110111101101101010100",
						 "100110111101101010011011",
						 "100110111101100111100010",
						 "100110111110010011001000",
						 "100110111110010000001110",
						 "100110111110001101010100",
						 "100110111110001010011010",
						 "100110111110000111100000",
						 "100110111110000100100110",
						 "100110111110000001101100",
						 "100110111101111110110010",
						 "100110111101111011111000",
						 "100110111101111000111110",
						 "100110111101110110000100",
						 "100110111101110011001010",
						 "100110111101110000010000",
						 "100110111101101101010110",
						 "100110111101101010011100",
						 "100110111101100111100010",
						 "100110111011110000001010",
						 "100110111011101101010000",
						 "100110111011101010010110",
						 "100110111011100111011100",
						 "100110111011100100100010",
						 "100110111011100001101000",
						 "100110111011011110101110",
						 "100110111011011011110100",
						 "100110111011011000111010",
						 "100110111011010110000000",
						 "100110111011010011000110",
						 "100110111011010000001100",
						 "100110111011001101010010",
						 "100110111011001010011000",
						 "100110111011000111011110",
						 "100110111011000100100100",
						 "100110111011110000001010",
						 "100110111011101101010000",
						 "100110111011101010010110",
						 "100110111011100111011100",
						 "100110111011100100100010",
						 "100110111011100001101000",
						 "100110111011011110101110",
						 "100110111011011011110100",
						 "100110111011011000111010",
						 "100110111011010110000000",
						 "100110111011010011000110",
						 "100110111011010000001100",
						 "100110111011001101010010",
						 "100110111011001010011000",
						 "100110111011000111011110",
						 "100110111011000100100100",
						 "100110111011110000001010",
						 "100110111011101101010000",
						 "100110111011101010010110",
						 "100110111011100111011100",
						 "100110111011100100100010",
						 "100110111011100001101000",
						 "100110111011011110101110",
						 "100110111011011011110100",
						 "100110111011011000111010",
						 "100110111011010110000000",
						 "100110111011010011000110",
						 "100110111011010000001100",
						 "100110111011001101010010",
						 "100110111011001010011000",
						 "100110111011000111011110",
						 "100110111011000100100100",
						 "100110111011110000011001",
						 "100110111011101101011110",
						 "100110111011101010100011",
						 "100110111011100111101000",
						 "100110111011100100101101",
						 "100110111011100001110010",
						 "100110111011011110110111",
						 "100110111011011011111100",
						 "100110111011011001000001",
						 "100110111011010110000110",
						 "100110111011010011001011",
						 "100110111011010000010000",
						 "100110111011001101010101",
						 "100110111011001010011010",
						 "100110111011000111011111",
						 "100110111011000100100100",
						 "100110111001001101011011",
						 "100110111001001010100000",
						 "100110111001000111100101",
						 "100110111001000100101010",
						 "100110111001000001101111",
						 "100110111000111110110100",
						 "100110111000111011111001",
						 "100110111000111000111110",
						 "100110111000110110000011",
						 "100110111000110011001000",
						 "100110111000110000001101",
						 "100110111000101101010010",
						 "100110111000101010010111",
						 "100110111000100111011100",
						 "100110111000100100100001",
						 "100110111000100001100110",
						 "100110111001001101011011",
						 "100110111001001010100000",
						 "100110111001000111100101",
						 "100110111001000100101010",
						 "100110111001000001101111",
						 "100110111000111110110100",
						 "100110111000111011111001",
						 "100110111000111000111110",
						 "100110111000110110000011",
						 "100110111000110011001000",
						 "100110111000110000001101",
						 "100110111000101101010010",
						 "100110111000101010010111",
						 "100110111000100111011100",
						 "100110111000100100100001",
						 "100110111000100001100110",
						 "100110111001001101011011",
						 "100110111001001010100000",
						 "100110111001000111100101",
						 "100110111001000100101010",
						 "100110111001000001101111",
						 "100110111000111110110100",
						 "100110111000111011111001",
						 "100110111000111000111110",
						 "100110111000110110000011",
						 "100110111000110011001000",
						 "100110111000110000001101",
						 "100110111000101101010010",
						 "100110111000101010010111",
						 "100110111000100111011100",
						 "100110111000100100100001",
						 "100110111000100001100110",
						 "100110110110101010101100",
						 "100110110110100111110000",
						 "100110110110100100110100",
						 "100110110110100001111000",
						 "100110110110011110111100",
						 "100110110110011100000000",
						 "100110110110011001000100",
						 "100110110110010110001000",
						 "100110110110010011001100",
						 "100110110110010000010000",
						 "100110110110001101010100",
						 "100110110110001010011000",
						 "100110110110000111011100",
						 "100110110110000100100000",
						 "100110110110000001100100",
						 "100110110101111110101000",
						 "100110110110101010101100",
						 "100110110110100111110000",
						 "100110110110100100110100",
						 "100110110110100001111000",
						 "100110110110011110111100",
						 "100110110110011100000000",
						 "100110110110011001000100",
						 "100110110110010110001000",
						 "100110110110010011001100",
						 "100110110110010000010000",
						 "100110110110001101010100",
						 "100110110110001010011000",
						 "100110110110000111011100",
						 "100110110110000100100000",
						 "100110110110000001100100",
						 "100110110101111110101000",
						 "100110110110101010101100",
						 "100110110110100111110000",
						 "100110110110100100110100",
						 "100110110110100001111000",
						 "100110110110011110111100",
						 "100110110110011100000000",
						 "100110110110011001000100",
						 "100110110110010110001000",
						 "100110110110010011001100",
						 "100110110110010000010000",
						 "100110110110001101010100",
						 "100110110110001010011000",
						 "100110110110000111011100",
						 "100110110110000100100000",
						 "100110110110000001100100",
						 "100110110101111110101000",
						 "100110110110101010111011",
						 "100110110110100111111110",
						 "100110110110100101000001",
						 "100110110110100010000100",
						 "100110110110011111000111",
						 "100110110110011100001010",
						 "100110110110011001001101",
						 "100110110110010110010000",
						 "100110110110010011010011",
						 "100110110110010000010110",
						 "100110110110001101011001",
						 "100110110110001010011100",
						 "100110110110000111011111",
						 "100110110110000100100010",
						 "100110110110000001100101",
						 "100110110101111110101000",
						 "100110110100000111111101",
						 "100110110100000101000000",
						 "100110110100000010000011",
						 "100110110011111111000110",
						 "100110110011111100001001",
						 "100110110011111001001100",
						 "100110110011110110001111",
						 "100110110011110011010010",
						 "100110110011110000010101",
						 "100110110011101101011000",
						 "100110110011101010011011",
						 "100110110011100111011110",
						 "100110110011100100100001",
						 "100110110011100001100100",
						 "100110110011011110100111",
						 "100110110011011011101010",
						 "100110110100000111111101",
						 "100110110100000101000000",
						 "100110110100000010000011",
						 "100110110011111111000110",
						 "100110110011111100001001",
						 "100110110011111001001100",
						 "100110110011110110001111",
						 "100110110011110011010010",
						 "100110110011110000010101",
						 "100110110011101101011000",
						 "100110110011101010011011",
						 "100110110011100111011110",
						 "100110110011100100100001",
						 "100110110011100001100100",
						 "100110110011011110100111",
						 "100110110011011011101010",
						 "100110110100000111111101",
						 "100110110100000101000000",
						 "100110110100000010000011",
						 "100110110011111111000110",
						 "100110110011111100001001",
						 "100110110011111001001100",
						 "100110110011110110001111",
						 "100110110011110011010010",
						 "100110110011110000010101",
						 "100110110011101101011000",
						 "100110110011101010011011",
						 "100110110011100111011110",
						 "100110110011100100100001",
						 "100110110011100001100100",
						 "100110110011011110100111",
						 "100110110011011011101010",
						 "100110110001100101001110",
						 "100110110001100010010000",
						 "100110110001011111010010",
						 "100110110001011100010100",
						 "100110110001011001010110",
						 "100110110001010110011000",
						 "100110110001010011011010",
						 "100110110001010000011100",
						 "100110110001001101011110",
						 "100110110001001010100000",
						 "100110110001000111100010",
						 "100110110001000100100100",
						 "100110110001000001100110",
						 "100110110000111110101000",
						 "100110110000111011101010",
						 "100110110000111000101100",
						 "100110110001100101001110",
						 "100110110001100010010000",
						 "100110110001011111010010",
						 "100110110001011100010100",
						 "100110110001011001010110",
						 "100110110001010110011000",
						 "100110110001010011011010",
						 "100110110001010000011100",
						 "100110110001001101011110",
						 "100110110001001010100000",
						 "100110110001000111100010",
						 "100110110001000100100100",
						 "100110110001000001100110",
						 "100110110000111110101000",
						 "100110110000111011101010",
						 "100110110000111000101100",
						 "100110110001100101001110",
						 "100110110001100010010000",
						 "100110110001011111010010",
						 "100110110001011100010100",
						 "100110110001011001010110",
						 "100110110001010110011000",
						 "100110110001010011011010",
						 "100110110001010000011100",
						 "100110110001001101011110",
						 "100110110001001010100000",
						 "100110110001000111100010",
						 "100110110001000100100100",
						 "100110110001000001100110",
						 "100110110000111110101000",
						 "100110110000111011101010",
						 "100110110000111000101100",
						 "100110110001100101001110",
						 "100110110001100010010000",
						 "100110110001011111010010",
						 "100110110001011100010100",
						 "100110110001011001010110",
						 "100110110001010110011000",
						 "100110110001010011011010",
						 "100110110001010000011100",
						 "100110110001001101011110",
						 "100110110001001010100000",
						 "100110110001000111100010",
						 "100110110001000100100100",
						 "100110110001000001100110",
						 "100110110000111110101000",
						 "100110110000111011101010",
						 "100110110000111000101100",
						 "100110101111000010011111",
						 "100110101110111111100000",
						 "100110101110111100100001",
						 "100110101110111001100010",
						 "100110101110110110100011",
						 "100110101110110011100100",
						 "100110101110110000100101",
						 "100110101110101101100110",
						 "100110101110101010100111",
						 "100110101110100111101000",
						 "100110101110100100101001",
						 "100110101110100001101010",
						 "100110101110011110101011",
						 "100110101110011011101100",
						 "100110101110011000101101",
						 "100110101110010101101110",
						 "100110101111000010011111",
						 "100110101110111111100000",
						 "100110101110111100100001",
						 "100110101110111001100010",
						 "100110101110110110100011",
						 "100110101110110011100100",
						 "100110101110110000100101",
						 "100110101110101101100110",
						 "100110101110101010100111",
						 "100110101110100111101000",
						 "100110101110100100101001",
						 "100110101110100001101010",
						 "100110101110011110101011",
						 "100110101110011011101100",
						 "100110101110011000101101",
						 "100110101110010101101110",
						 "100110101111000010011111",
						 "100110101110111111100000",
						 "100110101110111100100001",
						 "100110101110111001100010",
						 "100110101110110110100011",
						 "100110101110110011100100",
						 "100110101110110000100101",
						 "100110101110101101100110",
						 "100110101110101010100111",
						 "100110101110100111101000",
						 "100110101110100100101001",
						 "100110101110100001101010",
						 "100110101110011110101011",
						 "100110101110011011101100",
						 "100110101110011000101101",
						 "100110101110010101101110",
						 "100110101100011111100001",
						 "100110101100011100100010",
						 "100110101100011001100011",
						 "100110101100010110100100",
						 "100110101100010011100101",
						 "100110101100010000100110",
						 "100110101100001101100111",
						 "100110101100001010101000",
						 "100110101100000111101001",
						 "100110101100000100101010",
						 "100110101100000001101011",
						 "100110101011111110101100",
						 "100110101011111011101101",
						 "100110101011111000101110",
						 "100110101011110101101111",
						 "100110101011110010110000",
						 "100110101100011111110000",
						 "100110101100011100110000",
						 "100110101100011001110000",
						 "100110101100010110110000",
						 "100110101100010011110000",
						 "100110101100010000110000",
						 "100110101100001101110000",
						 "100110101100001010110000",
						 "100110101100000111110000",
						 "100110101100000100110000",
						 "100110101100000001110000",
						 "100110101011111110110000",
						 "100110101011111011110000",
						 "100110101011111000110000",
						 "100110101011110101110000",
						 "100110101011110010110000",
						 "100110101100011111110000",
						 "100110101100011100110000",
						 "100110101100011001110000",
						 "100110101100010110110000",
						 "100110101100010011110000",
						 "100110101100010000110000",
						 "100110101100001101110000",
						 "100110101100001010110000",
						 "100110101100000111110000",
						 "100110101100000100110000",
						 "100110101100000001110000",
						 "100110101011111110110000",
						 "100110101011111011110000",
						 "100110101011111000110000",
						 "100110101011110101110000",
						 "100110101011110010110000",
						 "100110101001111100110010",
						 "100110101001111001110010",
						 "100110101001110110110010",
						 "100110101001110011110010",
						 "100110101001110000110010",
						 "100110101001101101110010",
						 "100110101001101010110010",
						 "100110101001100111110010",
						 "100110101001100100110010",
						 "100110101001100001110010",
						 "100110101001011110110010",
						 "100110101001011011110010",
						 "100110101001011000110010",
						 "100110101001010101110010",
						 "100110101001010010110010",
						 "100110101001001111110010",
						 "100110101001111100110010",
						 "100110101001111001110010",
						 "100110101001110110110010",
						 "100110101001110011110010",
						 "100110101001110000110010",
						 "100110101001101101110010",
						 "100110101001101010110010",
						 "100110101001100111110010",
						 "100110101001100100110010",
						 "100110101001100001110010",
						 "100110101001011110110010",
						 "100110101001011011110010",
						 "100110101001011000110010",
						 "100110101001010101110010",
						 "100110101001010010110010",
						 "100110101001001111110010",
						 "100110101001111101000001",
						 "100110101001111010000000",
						 "100110101001110110111111",
						 "100110101001110011111110",
						 "100110101001110000111101",
						 "100110101001101101111100",
						 "100110101001101010111011",
						 "100110101001100111111010",
						 "100110101001100100111001",
						 "100110101001100001111000",
						 "100110101001011110110111",
						 "100110101001011011110110",
						 "100110101001011000110101",
						 "100110101001010101110100",
						 "100110101001010010110011",
						 "100110101001001111110010",
						 "100110101001111101000001",
						 "100110101001111010000000",
						 "100110101001110110111111",
						 "100110101001110011111110",
						 "100110101001110000111101",
						 "100110101001101101111100",
						 "100110101001101010111011",
						 "100110101001100111111010",
						 "100110101001100100111001",
						 "100110101001100001111000",
						 "100110101001011110110111",
						 "100110101001011011110110",
						 "100110101001011000110101",
						 "100110101001010101110100",
						 "100110101001010010110011",
						 "100110101001001111110010",
						 "100110100111011010000011",
						 "100110100111010111000010",
						 "100110100111010100000001",
						 "100110100111010001000000",
						 "100110100111001101111111",
						 "100110100111001010111110",
						 "100110100111000111111101",
						 "100110100111000100111100",
						 "100110100111000001111011",
						 "100110100110111110111010",
						 "100110100110111011111001",
						 "100110100110111000111000",
						 "100110100110110101110111",
						 "100110100110110010110110",
						 "100110100110101111110101",
						 "100110100110101100110100",
						 "100110100111011010000011",
						 "100110100111010111000010",
						 "100110100111010100000001",
						 "100110100111010001000000",
						 "100110100111001101111111",
						 "100110100111001010111110",
						 "100110100111000111111101",
						 "100110100111000100111100",
						 "100110100111000001111011",
						 "100110100110111110111010",
						 "100110100110111011111001",
						 "100110100110111000111000",
						 "100110100110110101110111",
						 "100110100110110010110110",
						 "100110100110101111110101",
						 "100110100110101100110100",
						 "100110100111011010010010",
						 "100110100111010111010000",
						 "100110100111010100001110",
						 "100110100111010001001100",
						 "100110100111001110001010",
						 "100110100111001011001000",
						 "100110100111001000000110",
						 "100110100111000101000100",
						 "100110100111000010000010",
						 "100110100110111111000000",
						 "100110100110111011111110",
						 "100110100110111000111100",
						 "100110100110110101111010",
						 "100110100110110010111000",
						 "100110100110101111110110",
						 "100110100110101100110100",
						 "100110100100110111010100",
						 "100110100100110100010010",
						 "100110100100110001010000",
						 "100110100100101110001110",
						 "100110100100101011001100",
						 "100110100100101000001010",
						 "100110100100100101001000",
						 "100110100100100010000110",
						 "100110100100011111000100",
						 "100110100100011100000010",
						 "100110100100011001000000",
						 "100110100100010101111110",
						 "100110100100010010111100",
						 "100110100100001111111010",
						 "100110100100001100111000",
						 "100110100100001001110110",
						 "100110100100110111010100",
						 "100110100100110100010010",
						 "100110100100110001010000",
						 "100110100100101110001110",
						 "100110100100101011001100",
						 "100110100100101000001010",
						 "100110100100100101001000",
						 "100110100100100010000110",
						 "100110100100011111000100",
						 "100110100100011100000010",
						 "100110100100011001000000",
						 "100110100100010101111110",
						 "100110100100010010111100",
						 "100110100100001111111010",
						 "100110100100001100111000",
						 "100110100100001001110110",
						 "100110100100110111010100",
						 "100110100100110100010010",
						 "100110100100110001010000",
						 "100110100100101110001110",
						 "100110100100101011001100",
						 "100110100100101000001010",
						 "100110100100100101001000",
						 "100110100100100010000110",
						 "100110100100011111000100",
						 "100110100100011100000010",
						 "100110100100011001000000",
						 "100110100100010101111110",
						 "100110100100010010111100",
						 "100110100100001111111010",
						 "100110100100001100111000",
						 "100110100100001001110110",
						 "100110100010010100100101",
						 "100110100010010001100010",
						 "100110100010001110011111",
						 "100110100010001011011100",
						 "100110100010001000011001",
						 "100110100010000101010110",
						 "100110100010000010010011",
						 "100110100001111111010000",
						 "100110100001111100001101",
						 "100110100001111001001010",
						 "100110100001110110000111",
						 "100110100001110011000100",
						 "100110100001110000000001",
						 "100110100001101100111110",
						 "100110100001101001111011",
						 "100110100001100110111000",
						 "100110100010010100100101",
						 "100110100010010001100010",
						 "100110100010001110011111",
						 "100110100010001011011100",
						 "100110100010001000011001",
						 "100110100010000101010110",
						 "100110100010000010010011",
						 "100110100001111111010000",
						 "100110100001111100001101",
						 "100110100001111001001010",
						 "100110100001110110000111",
						 "100110100001110011000100",
						 "100110100001110000000001",
						 "100110100001101100111110",
						 "100110100001101001111011",
						 "100110100001100110111000",
						 "100110100010010100100101",
						 "100110100010010001100010",
						 "100110100010001110011111",
						 "100110100010001011011100",
						 "100110100010001000011001",
						 "100110100010000101010110",
						 "100110100010000010010011",
						 "100110100001111111010000",
						 "100110100001111100001101",
						 "100110100001111001001010",
						 "100110100001110110000111",
						 "100110100001110011000100",
						 "100110100001110000000001",
						 "100110100001101100111110",
						 "100110100001101001111011",
						 "100110100001100110111000",
						 "100110100010010100100101",
						 "100110100010010001100010",
						 "100110100010001110011111",
						 "100110100010001011011100",
						 "100110100010001000011001",
						 "100110100010000101010110",
						 "100110100010000010010011",
						 "100110100001111111010000",
						 "100110100001111100001101",
						 "100110100001111001001010",
						 "100110100001110110000111",
						 "100110100001110011000100",
						 "100110100001110000000001",
						 "100110100001101100111110",
						 "100110100001101001111011",
						 "100110100001100110111000",
						 "100110011111110001110110",
						 "100110011111101110110010",
						 "100110011111101011101110",
						 "100110011111101000101010",
						 "100110011111100101100110",
						 "100110011111100010100010",
						 "100110011111011111011110",
						 "100110011111011100011010",
						 "100110011111011001010110",
						 "100110011111010110010010",
						 "100110011111010011001110",
						 "100110011111010000001010",
						 "100110011111001101000110",
						 "100110011111001010000010",
						 "100110011111000110111110",
						 "100110011111000011111010",
						 "100110011111110001110110",
						 "100110011111101110110010",
						 "100110011111101011101110",
						 "100110011111101000101010",
						 "100110011111100101100110",
						 "100110011111100010100010",
						 "100110011111011111011110",
						 "100110011111011100011010",
						 "100110011111011001010110",
						 "100110011111010110010010",
						 "100110011111010011001110",
						 "100110011111010000001010",
						 "100110011111001101000110",
						 "100110011111001010000010",
						 "100110011111000110111110",
						 "100110011111000011111010",
						 "100110011111110001110110",
						 "100110011111101110110010",
						 "100110011111101011101110",
						 "100110011111101000101010",
						 "100110011111100101100110",
						 "100110011111100010100010",
						 "100110011111011111011110",
						 "100110011111011100011010",
						 "100110011111011001010110",
						 "100110011111010110010010",
						 "100110011111010011001110",
						 "100110011111010000001010",
						 "100110011111001101000110",
						 "100110011111001010000010",
						 "100110011111000110111110",
						 "100110011111000011111010",
						 "100110011101001110111000",
						 "100110011101001011110100",
						 "100110011101001000110000",
						 "100110011101000101101100",
						 "100110011101000010101000",
						 "100110011100111111100100",
						 "100110011100111100100000",
						 "100110011100111001011100",
						 "100110011100110110011000",
						 "100110011100110011010100",
						 "100110011100110000010000",
						 "100110011100101101001100",
						 "100110011100101010001000",
						 "100110011100100111000100",
						 "100110011100100100000000",
						 "100110011100100000111100",
						 "100110011101001111000111",
						 "100110011101001100000010",
						 "100110011101001000111101",
						 "100110011101000101111000",
						 "100110011101000010110011",
						 "100110011100111111101110",
						 "100110011100111100101001",
						 "100110011100111001100100",
						 "100110011100110110011111",
						 "100110011100110011011010",
						 "100110011100110000010101",
						 "100110011100101101010000",
						 "100110011100101010001011",
						 "100110011100100111000110",
						 "100110011100100100000001",
						 "100110011100100000111100",
						 "100110011101001111000111",
						 "100110011101001100000010",
						 "100110011101001000111101",
						 "100110011101000101111000",
						 "100110011101000010110011",
						 "100110011100111111101110",
						 "100110011100111100101001",
						 "100110011100111001100100",
						 "100110011100110110011111",
						 "100110011100110011011010",
						 "100110011100110000010101",
						 "100110011100101101010000",
						 "100110011100101010001011",
						 "100110011100100111000110",
						 "100110011100100100000001",
						 "100110011100100000111100",
						 "100110011010101100001001",
						 "100110011010101001000100",
						 "100110011010100101111111",
						 "100110011010100010111010",
						 "100110011010011111110101",
						 "100110011010011100110000",
						 "100110011010011001101011",
						 "100110011010010110100110",
						 "100110011010010011100001",
						 "100110011010010000011100",
						 "100110011010001101010111",
						 "100110011010001010010010",
						 "100110011010000111001101",
						 "100110011010000100001000",
						 "100110011010000001000011",
						 "100110011001111101111110",
						 "100110011010101100001001",
						 "100110011010101001000100",
						 "100110011010100101111111",
						 "100110011010100010111010",
						 "100110011010011111110101",
						 "100110011010011100110000",
						 "100110011010011001101011",
						 "100110011010010110100110",
						 "100110011010010011100001",
						 "100110011010010000011100",
						 "100110011010001101010111",
						 "100110011010001010010010",
						 "100110011010000111001101",
						 "100110011010000100001000",
						 "100110011010000001000011",
						 "100110011001111101111110",
						 "100110011010101100011000",
						 "100110011010101001010010",
						 "100110011010100110001100",
						 "100110011010100011000110",
						 "100110011010100000000000",
						 "100110011010011100111010",
						 "100110011010011001110100",
						 "100110011010010110101110",
						 "100110011010010011101000",
						 "100110011010010000100010",
						 "100110011010001101011100",
						 "100110011010001010010110",
						 "100110011010000111010000",
						 "100110011010000100001010",
						 "100110011010000001000100",
						 "100110011001111101111110",
						 "100110011010101100011000",
						 "100110011010101001010010",
						 "100110011010100110001100",
						 "100110011010100011000110",
						 "100110011010100000000000",
						 "100110011010011100111010",
						 "100110011010011001110100",
						 "100110011010010110101110",
						 "100110011010010011101000",
						 "100110011010010000100010",
						 "100110011010001101011100",
						 "100110011010001010010110",
						 "100110011010000111010000",
						 "100110011010000100001010",
						 "100110011010000001000100",
						 "100110011001111101111110",
						 "100110011000001001011010",
						 "100110011000000110010100",
						 "100110011000000011001110",
						 "100110011000000000001000",
						 "100110010111111101000010",
						 "100110010111111001111100",
						 "100110010111110110110110",
						 "100110010111110011110000",
						 "100110010111110000101010",
						 "100110010111101101100100",
						 "100110010111101010011110",
						 "100110010111100111011000",
						 "100110010111100100010010",
						 "100110010111100001001100",
						 "100110010111011110000110",
						 "100110010111011011000000",
						 "100110011000001001011010",
						 "100110011000000110010100",
						 "100110011000000011001110",
						 "100110011000000000001000",
						 "100110010111111101000010",
						 "100110010111111001111100",
						 "100110010111110110110110",
						 "100110010111110011110000",
						 "100110010111110000101010",
						 "100110010111101101100100",
						 "100110010111101010011110",
						 "100110010111100111011000",
						 "100110010111100100010010",
						 "100110010111100001001100",
						 "100110010111011110000110",
						 "100110010111011011000000",
						 "100110011000001001101001",
						 "100110011000000110100010",
						 "100110011000000011011011",
						 "100110011000000000010100",
						 "100110010111111101001101",
						 "100110010111111010000110",
						 "100110010111110110111111",
						 "100110010111110011111000",
						 "100110010111110000110001",
						 "100110010111101101101010",
						 "100110010111101010100011",
						 "100110010111100111011100",
						 "100110010111100100010101",
						 "100110010111100001001110",
						 "100110010111011110000111",
						 "100110010111011011000000",
						 "100110010101100110101011",
						 "100110010101100011100100",
						 "100110010101100000011101",
						 "100110010101011101010110",
						 "100110010101011010001111",
						 "100110010101010111001000",
						 "100110010101010100000001",
						 "100110010101010000111010",
						 "100110010101001101110011",
						 "100110010101001010101100",
						 "100110010101000111100101",
						 "100110010101000100011110",
						 "100110010101000001010111",
						 "100110010100111110010000",
						 "100110010100111011001001",
						 "100110010100111000000010",
						 "100110010101100110101011",
						 "100110010101100011100100",
						 "100110010101100000011101",
						 "100110010101011101010110",
						 "100110010101011010001111",
						 "100110010101010111001000",
						 "100110010101010100000001",
						 "100110010101010000111010",
						 "100110010101001101110011",
						 "100110010101001010101100",
						 "100110010101000111100101",
						 "100110010101000100011110",
						 "100110010101000001010111",
						 "100110010100111110010000",
						 "100110010100111011001001",
						 "100110010100111000000010",
						 "100110010101100110101011",
						 "100110010101100011100100",
						 "100110010101100000011101",
						 "100110010101011101010110",
						 "100110010101011010001111",
						 "100110010101010111001000",
						 "100110010101010100000001",
						 "100110010101010000111010",
						 "100110010101001101110011",
						 "100110010101001010101100",
						 "100110010101000111100101",
						 "100110010101000100011110",
						 "100110010101000001010111",
						 "100110010100111110010000",
						 "100110010100111011001001",
						 "100110010100111000000010",
						 "100110010011000011111100",
						 "100110010011000000110100",
						 "100110010010111101101100",
						 "100110010010111010100100",
						 "100110010010110111011100",
						 "100110010010110100010100",
						 "100110010010110001001100",
						 "100110010010101110000100",
						 "100110010010101010111100",
						 "100110010010100111110100",
						 "100110010010100100101100",
						 "100110010010100001100100",
						 "100110010010011110011100",
						 "100110010010011011010100",
						 "100110010010011000001100",
						 "100110010010010101000100",
						 "100110010011000011111100",
						 "100110010011000000110100",
						 "100110010010111101101100",
						 "100110010010111010100100",
						 "100110010010110111011100",
						 "100110010010110100010100",
						 "100110010010110001001100",
						 "100110010010101110000100",
						 "100110010010101010111100",
						 "100110010010100111110100",
						 "100110010010100100101100",
						 "100110010010100001100100",
						 "100110010010011110011100",
						 "100110010010011011010100",
						 "100110010010011000001100",
						 "100110010010010101000100",
						 "100110010011000011111100",
						 "100110010011000000110100",
						 "100110010010111101101100",
						 "100110010010111010100100",
						 "100110010010110111011100",
						 "100110010010110100010100",
						 "100110010010110001001100",
						 "100110010010101110000100",
						 "100110010010101010111100",
						 "100110010010100111110100",
						 "100110010010100100101100",
						 "100110010010100001100100",
						 "100110010010011110011100",
						 "100110010010011011010100",
						 "100110010010011000001100",
						 "100110010010010101000100",
						 "100110010011000011111100",
						 "100110010011000000110100",
						 "100110010010111101101100",
						 "100110010010111010100100",
						 "100110010010110111011100",
						 "100110010010110100010100",
						 "100110010010110001001100",
						 "100110010010101110000100",
						 "100110010010101010111100",
						 "100110010010100111110100",
						 "100110010010100100101100",
						 "100110010010100001100100",
						 "100110010010011110011100",
						 "100110010010011011010100",
						 "100110010010011000001100",
						 "100110010010010101000100",
						 "100110010000100001001101",
						 "100110010000011110000100",
						 "100110010000011010111011",
						 "100110010000010111110010",
						 "100110010000010100101001",
						 "100110010000010001100000",
						 "100110010000001110010111",
						 "100110010000001011001110",
						 "100110010000001000000101",
						 "100110010000000100111100",
						 "100110010000000001110011",
						 "100110001111111110101010",
						 "100110001111111011100001",
						 "100110001111111000011000",
						 "100110001111110101001111",
						 "100110001111110010000110",
						 "100110010000100001001101",
						 "100110010000011110000100",
						 "100110010000011010111011",
						 "100110010000010111110010",
						 "100110010000010100101001",
						 "100110010000010001100000",
						 "100110010000001110010111",
						 "100110010000001011001110",
						 "100110010000001000000101",
						 "100110010000000100111100",
						 "100110010000000001110011",
						 "100110001111111110101010",
						 "100110001111111011100001",
						 "100110001111111000011000",
						 "100110001111110101001111",
						 "100110001111110010000110",
						 "100110010000100001001101",
						 "100110010000011110000100",
						 "100110010000011010111011",
						 "100110010000010111110010",
						 "100110010000010100101001",
						 "100110010000010001100000",
						 "100110010000001110010111",
						 "100110010000001011001110",
						 "100110010000001000000101",
						 "100110010000000100111100",
						 "100110010000000001110011",
						 "100110001111111110101010",
						 "100110001111111011100001",
						 "100110001111111000011000",
						 "100110001111110101001111",
						 "100110001111110010000110",
						 "100110001101111110001111",
						 "100110001101111011000110",
						 "100110001101110111111101",
						 "100110001101110100110100",
						 "100110001101110001101011",
						 "100110001101101110100010",
						 "100110001101101011011001",
						 "100110001101101000010000",
						 "100110001101100101000111",
						 "100110001101100001111110",
						 "100110001101011110110101",
						 "100110001101011011101100",
						 "100110001101011000100011",
						 "100110001101010101011010",
						 "100110001101010010010001",
						 "100110001101001111001000",
						 "100110001101111110011110",
						 "100110001101111011010100",
						 "100110001101111000001010",
						 "100110001101110101000000",
						 "100110001101110001110110",
						 "100110001101101110101100",
						 "100110001101101011100010",
						 "100110001101101000011000",
						 "100110001101100101001110",
						 "100110001101100010000100",
						 "100110001101011110111010",
						 "100110001101011011110000",
						 "100110001101011000100110",
						 "100110001101010101011100",
						 "100110001101010010010010",
						 "100110001101001111001000",
						 "100110001101111110011110",
						 "100110001101111011010100",
						 "100110001101111000001010",
						 "100110001101110101000000",
						 "100110001101110001110110",
						 "100110001101101110101100",
						 "100110001101101011100010",
						 "100110001101101000011000",
						 "100110001101100101001110",
						 "100110001101100010000100",
						 "100110001101011110111010",
						 "100110001101011011110000",
						 "100110001101011000100110",
						 "100110001101010101011100",
						 "100110001101010010010010",
						 "100110001101001111001000",
						 "100110001011011011100000",
						 "100110001011011000010110",
						 "100110001011010101001100",
						 "100110001011010010000010",
						 "100110001011001110111000",
						 "100110001011001011101110",
						 "100110001011001000100100",
						 "100110001011000101011010",
						 "100110001011000010010000",
						 "100110001010111111000110",
						 "100110001010111011111100",
						 "100110001010111000110010",
						 "100110001010110101101000",
						 "100110001010110010011110",
						 "100110001010101111010100",
						 "100110001010101100001010",
						 "100110001011011011100000",
						 "100110001011011000010110",
						 "100110001011010101001100",
						 "100110001011010010000010",
						 "100110001011001110111000",
						 "100110001011001011101110",
						 "100110001011001000100100",
						 "100110001011000101011010",
						 "100110001011000010010000",
						 "100110001010111111000110",
						 "100110001010111011111100",
						 "100110001010111000110010",
						 "100110001010110101101000",
						 "100110001010110010011110",
						 "100110001010101111010100",
						 "100110001010101100001010",
						 "100110001011011011101111",
						 "100110001011011000100100",
						 "100110001011010101011001",
						 "100110001011010010001110",
						 "100110001011001111000011",
						 "100110001011001011111000",
						 "100110001011001000101101",
						 "100110001011000101100010",
						 "100110001011000010010111",
						 "100110001010111111001100",
						 "100110001010111100000001",
						 "100110001010111000110110",
						 "100110001010110101101011",
						 "100110001010110010100000",
						 "100110001010101111010101",
						 "100110001010101100001010",
						 "100110001000111000110001",
						 "100110001000110101100110",
						 "100110001000110010011011",
						 "100110001000101111010000",
						 "100110001000101100000101",
						 "100110001000101000111010",
						 "100110001000100101101111",
						 "100110001000100010100100",
						 "100110001000011111011001",
						 "100110001000011100001110",
						 "100110001000011001000011",
						 "100110001000010101111000",
						 "100110001000010010101101",
						 "100110001000001111100010",
						 "100110001000001100010111",
						 "100110001000001001001100",
						 "100110001000111000110001",
						 "100110001000110101100110",
						 "100110001000110010011011",
						 "100110001000101111010000",
						 "100110001000101100000101",
						 "100110001000101000111010",
						 "100110001000100101101111",
						 "100110001000100010100100",
						 "100110001000011111011001",
						 "100110001000011100001110",
						 "100110001000011001000011",
						 "100110001000010101111000",
						 "100110001000010010101101",
						 "100110001000001111100010",
						 "100110001000001100010111",
						 "100110001000001001001100",
						 "100110001000111000110001",
						 "100110001000110101100110",
						 "100110001000110010011011",
						 "100110001000101111010000",
						 "100110001000101100000101",
						 "100110001000101000111010",
						 "100110001000100101101111",
						 "100110001000100010100100",
						 "100110001000011111011001",
						 "100110001000011100001110",
						 "100110001000011001000011",
						 "100110001000010101111000",
						 "100110001000010010101101",
						 "100110001000001111100010",
						 "100110001000001100010111",
						 "100110001000001001001100",
						 "100110000110010110000010",
						 "100110000110010010110110",
						 "100110000110001111101010",
						 "100110000110001100011110",
						 "100110000110001001010010",
						 "100110000110000110000110",
						 "100110000110000010111010",
						 "100110000101111111101110",
						 "100110000101111100100010",
						 "100110000101111001010110",
						 "100110000101110110001010",
						 "100110000101110010111110",
						 "100110000101101111110010",
						 "100110000101101100100110",
						 "100110000101101001011010",
						 "100110000101100110001110",
						 "100110000110010110000010",
						 "100110000110010010110110",
						 "100110000110001111101010",
						 "100110000110001100011110",
						 "100110000110001001010010",
						 "100110000110000110000110",
						 "100110000110000010111010",
						 "100110000101111111101110",
						 "100110000101111100100010",
						 "100110000101111001010110",
						 "100110000101110110001010",
						 "100110000101110010111110",
						 "100110000101101111110010",
						 "100110000101101100100110",
						 "100110000101101001011010",
						 "100110000101100110001110",
						 "100110000110010110000010",
						 "100110000110010010110110",
						 "100110000110001111101010",
						 "100110000110001100011110",
						 "100110000110001001010010",
						 "100110000110000110000110",
						 "100110000110000010111010",
						 "100110000101111111101110",
						 "100110000101111100100010",
						 "100110000101111001010110",
						 "100110000101110110001010",
						 "100110000101110010111110",
						 "100110000101101111110010",
						 "100110000101101100100110",
						 "100110000101101001011010",
						 "100110000101100110001110",
						 "100110000110010110000010",
						 "100110000110010010110110",
						 "100110000110001111101010",
						 "100110000110001100011110",
						 "100110000110001001010010",
						 "100110000110000110000110",
						 "100110000110000010111010",
						 "100110000101111111101110",
						 "100110000101111100100010",
						 "100110000101111001010110",
						 "100110000101110110001010",
						 "100110000101110010111110",
						 "100110000101101111110010",
						 "100110000101101100100110",
						 "100110000101101001011010",
						 "100110000101100110001110",
						 "100110000011110011000100",
						 "100110000011101111111000",
						 "100110000011101100101100",
						 "100110000011101001100000",
						 "100110000011100110010100",
						 "100110000011100011001000",
						 "100110000011011111111100",
						 "100110000011011100110000",
						 "100110000011011001100100",
						 "100110000011010110011000",
						 "100110000011010011001100",
						 "100110000011010000000000",
						 "100110000011001100110100",
						 "100110000011001001101000",
						 "100110000011000110011100",
						 "100110000011000011010000",
						 "100110000011110011010011",
						 "100110000011110000000110",
						 "100110000011101100111001",
						 "100110000011101001101100",
						 "100110000011100110011111",
						 "100110000011100011010010",
						 "100110000011100000000101",
						 "100110000011011100111000",
						 "100110000011011001101011",
						 "100110000011010110011110",
						 "100110000011010011010001",
						 "100110000011010000000100",
						 "100110000011001100110111",
						 "100110000011001001101010",
						 "100110000011000110011101",
						 "100110000011000011010000",
						 "100110000011110011010011",
						 "100110000011110000000110",
						 "100110000011101100111001",
						 "100110000011101001101100",
						 "100110000011100110011111",
						 "100110000011100011010010",
						 "100110000011100000000101",
						 "100110000011011100111000",
						 "100110000011011001101011",
						 "100110000011010110011110",
						 "100110000011010011010001",
						 "100110000011010000000100",
						 "100110000011001100110111",
						 "100110000011001001101010",
						 "100110000011000110011101",
						 "100110000011000011010000",
						 "100110000001010000010101",
						 "100110000001001101001000",
						 "100110000001001001111011",
						 "100110000001000110101110",
						 "100110000001000011100001",
						 "100110000001000000010100",
						 "100110000000111101000111",
						 "100110000000111001111010",
						 "100110000000110110101101",
						 "100110000000110011100000",
						 "100110000000110000010011",
						 "100110000000101101000110",
						 "100110000000101001111001",
						 "100110000000100110101100",
						 "100110000000100011011111",
						 "100110000000100000010010",
						 "100110000001010000010101",
						 "100110000001001101001000",
						 "100110000001001001111011",
						 "100110000001000110101110",
						 "100110000001000011100001",
						 "100110000001000000010100",
						 "100110000000111101000111",
						 "100110000000111001111010",
						 "100110000000110110101101",
						 "100110000000110011100000",
						 "100110000000110000010011",
						 "100110000000101101000110",
						 "100110000000101001111001",
						 "100110000000100110101100",
						 "100110000000100011011111",
						 "100110000000100000010010",
						 "100110000001010000100100",
						 "100110000001001101010110",
						 "100110000001001010001000",
						 "100110000001000110111010",
						 "100110000001000011101100",
						 "100110000001000000011110",
						 "100110000000111101010000",
						 "100110000000111010000010",
						 "100110000000110110110100",
						 "100110000000110011100110",
						 "100110000000110000011000",
						 "100110000000101101001010",
						 "100110000000101001111100",
						 "100110000000100110101110",
						 "100110000000100011100000",
						 "100110000000100000010010",
						 "100101111110101101100110",
						 "100101111110101010011000",
						 "100101111110100111001010",
						 "100101111110100011111100",
						 "100101111110100000101110",
						 "100101111110011101100000",
						 "100101111110011010010010",
						 "100101111110010111000100",
						 "100101111110010011110110",
						 "100101111110010000101000",
						 "100101111110001101011010",
						 "100101111110001010001100",
						 "100101111110000110111110",
						 "100101111110000011110000",
						 "100101111110000000100010",
						 "100101111101111101010100",
						 "100101111110101101100110",
						 "100101111110101010011000",
						 "100101111110100111001010",
						 "100101111110100011111100",
						 "100101111110100000101110",
						 "100101111110011101100000",
						 "100101111110011010010010",
						 "100101111110010111000100",
						 "100101111110010011110110",
						 "100101111110010000101000",
						 "100101111110001101011010",
						 "100101111110001010001100",
						 "100101111110000110111110",
						 "100101111110000011110000",
						 "100101111110000000100010",
						 "100101111101111101010100",
						 "100101111110101101100110",
						 "100101111110101010011000",
						 "100101111110100111001010",
						 "100101111110100011111100",
						 "100101111110100000101110",
						 "100101111110011101100000",
						 "100101111110011010010010",
						 "100101111110010111000100",
						 "100101111110010011110110",
						 "100101111110010000101000",
						 "100101111110001101011010",
						 "100101111110001010001100",
						 "100101111110000110111110",
						 "100101111110000011110000",
						 "100101111110000000100010",
						 "100101111101111101010100",
						 "100101111100001010110111",
						 "100101111100000111101000",
						 "100101111100000100011001",
						 "100101111100000001001010",
						 "100101111011111101111011",
						 "100101111011111010101100",
						 "100101111011110111011101",
						 "100101111011110100001110",
						 "100101111011110000111111",
						 "100101111011101101110000",
						 "100101111011101010100001",
						 "100101111011100111010010",
						 "100101111011100100000011",
						 "100101111011100000110100",
						 "100101111011011101100101",
						 "100101111011011010010110",
						 "100101111100001010110111",
						 "100101111100000111101000",
						 "100101111100000100011001",
						 "100101111100000001001010",
						 "100101111011111101111011",
						 "100101111011111010101100",
						 "100101111011110111011101",
						 "100101111011110100001110",
						 "100101111011110000111111",
						 "100101111011101101110000",
						 "100101111011101010100001",
						 "100101111011100111010010",
						 "100101111011100100000011",
						 "100101111011100000110100",
						 "100101111011011101100101",
						 "100101111011011010010110",
						 "100101111100001010110111",
						 "100101111100000111101000",
						 "100101111100000100011001",
						 "100101111100000001001010",
						 "100101111011111101111011",
						 "100101111011111010101100",
						 "100101111011110111011101",
						 "100101111011110100001110",
						 "100101111011110000111111",
						 "100101111011101101110000",
						 "100101111011101010100001",
						 "100101111011100111010010",
						 "100101111011100100000011",
						 "100101111011100000110100",
						 "100101111011011101100101",
						 "100101111011011010010110",
						 "100101111001100111111001",
						 "100101111001100100101010",
						 "100101111001100001011011",
						 "100101111001011110001100",
						 "100101111001011010111101",
						 "100101111001010111101110",
						 "100101111001010100011111",
						 "100101111001010001010000",
						 "100101111001001110000001",
						 "100101111001001010110010",
						 "100101111001000111100011",
						 "100101111001000100010100",
						 "100101111001000001000101",
						 "100101111000111101110110",
						 "100101111000111010100111",
						 "100101111000110111011000",
						 "100101111001100111111001",
						 "100101111001100100101010",
						 "100101111001100001011011",
						 "100101111001011110001100",
						 "100101111001011010111101",
						 "100101111001010111101110",
						 "100101111001010100011111",
						 "100101111001010001010000",
						 "100101111001001110000001",
						 "100101111001001010110010",
						 "100101111001000111100011",
						 "100101111001000100010100",
						 "100101111001000001000101",
						 "100101111000111101110110",
						 "100101111000111010100111",
						 "100101111000110111011000",
						 "100101111001101000001000",
						 "100101111001100100111000",
						 "100101111001100001101000",
						 "100101111001011110011000",
						 "100101111001011011001000",
						 "100101111001010111111000",
						 "100101111001010100101000",
						 "100101111001010001011000",
						 "100101111001001110001000",
						 "100101111001001010111000",
						 "100101111001000111101000",
						 "100101111001000100011000",
						 "100101111001000001001000",
						 "100101111000111101111000",
						 "100101111000111010101000",
						 "100101111000110111011000",
						 "100101110111000101001010",
						 "100101110111000001111010",
						 "100101110110111110101010",
						 "100101110110111011011010",
						 "100101110110111000001010",
						 "100101110110110100111010",
						 "100101110110110001101010",
						 "100101110110101110011010",
						 "100101110110101011001010",
						 "100101110110100111111010",
						 "100101110110100100101010",
						 "100101110110100001011010",
						 "100101110110011110001010",
						 "100101110110011010111010",
						 "100101110110010111101010",
						 "100101110110010100011010",
						 "100101110111000101001010",
						 "100101110111000001111010",
						 "100101110110111110101010",
						 "100101110110111011011010",
						 "100101110110111000001010",
						 "100101110110110100111010",
						 "100101110110110001101010",
						 "100101110110101110011010",
						 "100101110110101011001010",
						 "100101110110100111111010",
						 "100101110110100100101010",
						 "100101110110100001011010",
						 "100101110110011110001010",
						 "100101110110011010111010",
						 "100101110110010111101010",
						 "100101110110010100011010",
						 "100101110111000101001010",
						 "100101110111000001111010",
						 "100101110110111110101010",
						 "100101110110111011011010",
						 "100101110110111000001010",
						 "100101110110110100111010",
						 "100101110110110001101010",
						 "100101110110101110011010",
						 "100101110110101011001010",
						 "100101110110100111111010",
						 "100101110110100100101010",
						 "100101110110100001011010",
						 "100101110110011110001010",
						 "100101110110011010111010",
						 "100101110110010111101010",
						 "100101110110010100011010",
						 "100101110111000101011001",
						 "100101110111000010001000",
						 "100101110110111110110111",
						 "100101110110111011100110",
						 "100101110110111000010101",
						 "100101110110110101000100",
						 "100101110110110001110011",
						 "100101110110101110100010",
						 "100101110110101011010001",
						 "100101110110101000000000",
						 "100101110110100100101111",
						 "100101110110100001011110",
						 "100101110110011110001101",
						 "100101110110011010111100",
						 "100101110110010111101011",
						 "100101110110010100011010",
						 "100101110100100010011011",
						 "100101110100011111001010",
						 "100101110100011011111001",
						 "100101110100011000101000",
						 "100101110100010101010111",
						 "100101110100010010000110",
						 "100101110100001110110101",
						 "100101110100001011100100",
						 "100101110100001000010011",
						 "100101110100000101000010",
						 "100101110100000001110001",
						 "100101110011111110100000",
						 "100101110011111011001111",
						 "100101110011110111111110",
						 "100101110011110100101101",
						 "100101110011110001011100",
						 "100101110100100010011011",
						 "100101110100011111001010",
						 "100101110100011011111001",
						 "100101110100011000101000",
						 "100101110100010101010111",
						 "100101110100010010000110",
						 "100101110100001110110101",
						 "100101110100001011100100",
						 "100101110100001000010011",
						 "100101110100000101000010",
						 "100101110100000001110001",
						 "100101110011111110100000",
						 "100101110011111011001111",
						 "100101110011110111111110",
						 "100101110011110100101101",
						 "100101110011110001011100",
						 "100101110100100010011011",
						 "100101110100011111001010",
						 "100101110100011011111001",
						 "100101110100011000101000",
						 "100101110100010101010111",
						 "100101110100010010000110",
						 "100101110100001110110101",
						 "100101110100001011100100",
						 "100101110100001000010011",
						 "100101110100000101000010",
						 "100101110100000001110001",
						 "100101110011111110100000",
						 "100101110011111011001111",
						 "100101110011110111111110",
						 "100101110011110100101101",
						 "100101110011110001011100",
						 "100101110001111111011101",
						 "100101110001111100001100",
						 "100101110001111000111011",
						 "100101110001110101101010",
						 "100101110001110010011001",
						 "100101110001101111001000",
						 "100101110001101011110111",
						 "100101110001101000100110",
						 "100101110001100101010101",
						 "100101110001100010000100",
						 "100101110001011110110011",
						 "100101110001011011100010",
						 "100101110001011000010001",
						 "100101110001010101000000",
						 "100101110001010001101111",
						 "100101110001001110011110",
						 "100101110001111111101100",
						 "100101110001111100011010",
						 "100101110001111001001000",
						 "100101110001110101110110",
						 "100101110001110010100100",
						 "100101110001101111010010",
						 "100101110001101100000000",
						 "100101110001101000101110",
						 "100101110001100101011100",
						 "100101110001100010001010",
						 "100101110001011110111000",
						 "100101110001011011100110",
						 "100101110001011000010100",
						 "100101110001010101000010",
						 "100101110001010001110000",
						 "100101110001001110011110",
						 "100101110001111111101100",
						 "100101110001111100011010",
						 "100101110001111001001000",
						 "100101110001110101110110",
						 "100101110001110010100100",
						 "100101110001101111010010",
						 "100101110001101100000000",
						 "100101110001101000101110",
						 "100101110001100101011100",
						 "100101110001100010001010",
						 "100101110001011110111000",
						 "100101110001011011100110",
						 "100101110001011000010100",
						 "100101110001010101000010",
						 "100101110001010001110000",
						 "100101110001001110011110",
						 "100101101111011100101110",
						 "100101101111011001011100",
						 "100101101111010110001010",
						 "100101101111010010111000",
						 "100101101111001111100110",
						 "100101101111001100010100",
						 "100101101111001001000010",
						 "100101101111000101110000",
						 "100101101111000010011110",
						 "100101101110111111001100",
						 "100101101110111011111010",
						 "100101101110111000101000",
						 "100101101110110101010110",
						 "100101101110110010000100",
						 "100101101110101110110010",
						 "100101101110101011100000",
						 "100101101111011100101110",
						 "100101101111011001011100",
						 "100101101111010110001010",
						 "100101101111010010111000",
						 "100101101111001111100110",
						 "100101101111001100010100",
						 "100101101111001001000010",
						 "100101101111000101110000",
						 "100101101111000010011110",
						 "100101101110111111001100",
						 "100101101110111011111010",
						 "100101101110111000101000",
						 "100101101110110101010110",
						 "100101101110110010000100",
						 "100101101110101110110010",
						 "100101101110101011100000",
						 "100101101111011100111101",
						 "100101101111011001101010",
						 "100101101111010110010111",
						 "100101101111010011000100",
						 "100101101111001111110001",
						 "100101101111001100011110",
						 "100101101111001001001011",
						 "100101101111000101111000",
						 "100101101111000010100101",
						 "100101101110111111010010",
						 "100101101110111011111111",
						 "100101101110111000101100",
						 "100101101110110101011001",
						 "100101101110110010000110",
						 "100101101110101110110011",
						 "100101101110101011100000",
						 "100101101100111001111111",
						 "100101101100110110101100",
						 "100101101100110011011001",
						 "100101101100110000000110",
						 "100101101100101100110011",
						 "100101101100101001100000",
						 "100101101100100110001101",
						 "100101101100100010111010",
						 "100101101100011111100111",
						 "100101101100011100010100",
						 "100101101100011001000001",
						 "100101101100010101101110",
						 "100101101100010010011011",
						 "100101101100001111001000",
						 "100101101100001011110101",
						 "100101101100001000100010",
						 "100101101100111001111111",
						 "100101101100110110101100",
						 "100101101100110011011001",
						 "100101101100110000000110",
						 "100101101100101100110011",
						 "100101101100101001100000",
						 "100101101100100110001101",
						 "100101101100100010111010",
						 "100101101100011111100111",
						 "100101101100011100010100",
						 "100101101100011001000001",
						 "100101101100010101101110",
						 "100101101100010010011011",
						 "100101101100001111001000",
						 "100101101100001011110101",
						 "100101101100001000100010",
						 "100101101100111001111111",
						 "100101101100110110101100",
						 "100101101100110011011001",
						 "100101101100110000000110",
						 "100101101100101100110011",
						 "100101101100101001100000",
						 "100101101100100110001101",
						 "100101101100100010111010",
						 "100101101100011111100111",
						 "100101101100011100010100",
						 "100101101100011001000001",
						 "100101101100010101101110",
						 "100101101100010010011011",
						 "100101101100001111001000",
						 "100101101100001011110101",
						 "100101101100001000100010",
						 "100101101010010111000001",
						 "100101101010010011101110",
						 "100101101010010000011011",
						 "100101101010001101001000",
						 "100101101010001001110101",
						 "100101101010000110100010",
						 "100101101010000011001111",
						 "100101101001111111111100",
						 "100101101001111100101001",
						 "100101101001111001010110",
						 "100101101001110110000011",
						 "100101101001110010110000",
						 "100101101001101111011101",
						 "100101101001101100001010",
						 "100101101001101000110111",
						 "100101101001100101100100",
						 "100101101010010111010000",
						 "100101101010010011111100",
						 "100101101010010000101000",
						 "100101101010001101010100",
						 "100101101010001010000000",
						 "100101101010000110101100",
						 "100101101010000011011000",
						 "100101101010000000000100",
						 "100101101001111100110000",
						 "100101101001111001011100",
						 "100101101001110110001000",
						 "100101101001110010110100",
						 "100101101001101111100000",
						 "100101101001101100001100",
						 "100101101001101000111000",
						 "100101101001100101100100",
						 "100101101010010111010000",
						 "100101101010010011111100",
						 "100101101010010000101000",
						 "100101101010001101010100",
						 "100101101010001010000000",
						 "100101101010000110101100",
						 "100101101010000011011000",
						 "100101101010000000000100",
						 "100101101001111100110000",
						 "100101101001111001011100",
						 "100101101001110110001000",
						 "100101101001110010110100",
						 "100101101001101111100000",
						 "100101101001101100001100",
						 "100101101001101000111000",
						 "100101101001100101100100",
						 "100101100111110100010010",
						 "100101100111110000111110",
						 "100101100111101101101010",
						 "100101100111101010010110",
						 "100101100111100111000010",
						 "100101100111100011101110",
						 "100101100111100000011010",
						 "100101100111011101000110",
						 "100101100111011001110010",
						 "100101100111010110011110",
						 "100101100111010011001010",
						 "100101100111001111110110",
						 "100101100111001100100010",
						 "100101100111001001001110",
						 "100101100111000101111010",
						 "100101100111000010100110",
						 "100101100111110100010010",
						 "100101100111110000111110",
						 "100101100111101101101010",
						 "100101100111101010010110",
						 "100101100111100111000010",
						 "100101100111100011101110",
						 "100101100111100000011010",
						 "100101100111011101000110",
						 "100101100111011001110010",
						 "100101100111010110011110",
						 "100101100111010011001010",
						 "100101100111001111110110",
						 "100101100111001100100010",
						 "100101100111001001001110",
						 "100101100111000101111010",
						 "100101100111000010100110",
						 "100101100111110100100001",
						 "100101100111110001001100",
						 "100101100111101101110111",
						 "100101100111101010100010",
						 "100101100111100111001101",
						 "100101100111100011111000",
						 "100101100111100000100011",
						 "100101100111011101001110",
						 "100101100111011001111001",
						 "100101100111010110100100",
						 "100101100111010011001111",
						 "100101100111001111111010",
						 "100101100111001100100101",
						 "100101100111001001010000",
						 "100101100111000101111011",
						 "100101100111000010100110",
						 "100101100101010001100011",
						 "100101100101001110001110",
						 "100101100101001010111001",
						 "100101100101000111100100",
						 "100101100101000100001111",
						 "100101100101000000111010",
						 "100101100100111101100101",
						 "100101100100111010010000",
						 "100101100100110110111011",
						 "100101100100110011100110",
						 "100101100100110000010001",
						 "100101100100101100111100",
						 "100101100100101001100111",
						 "100101100100100110010010",
						 "100101100100100010111101",
						 "100101100100011111101000",
						 "100101100101010001100011",
						 "100101100101001110001110",
						 "100101100101001010111001",
						 "100101100101000111100100",
						 "100101100101000100001111",
						 "100101100101000000111010",
						 "100101100100111101100101",
						 "100101100100111010010000",
						 "100101100100110110111011",
						 "100101100100110011100110",
						 "100101100100110000010001",
						 "100101100100101100111100",
						 "100101100100101001100111",
						 "100101100100100110010010",
						 "100101100100100010111101",
						 "100101100100011111101000",
						 "100101100101010001100011",
						 "100101100101001110001110",
						 "100101100101001010111001",
						 "100101100101000111100100",
						 "100101100101000100001111",
						 "100101100101000000111010",
						 "100101100100111101100101",
						 "100101100100111010010000",
						 "100101100100110110111011",
						 "100101100100110011100110",
						 "100101100100110000010001",
						 "100101100100101100111100",
						 "100101100100101001100111",
						 "100101100100100110010010",
						 "100101100100100010111101",
						 "100101100100011111101000",
						 "100101100010101110100101",
						 "100101100010101011010000",
						 "100101100010100111111011",
						 "100101100010100100100110",
						 "100101100010100001010001",
						 "100101100010011101111100",
						 "100101100010011010100111",
						 "100101100010010111010010",
						 "100101100010010011111101",
						 "100101100010010000101000",
						 "100101100010001101010011",
						 "100101100010001001111110",
						 "100101100010000110101001",
						 "100101100010000011010100",
						 "100101100001111111111111",
						 "100101100001111100101010",
						 "100101100010101110110100",
						 "100101100010101011011110",
						 "100101100010101000001000",
						 "100101100010100100110010",
						 "100101100010100001011100",
						 "100101100010011110000110",
						 "100101100010011010110000",
						 "100101100010010111011010",
						 "100101100010010100000100",
						 "100101100010010000101110",
						 "100101100010001101011000",
						 "100101100010001010000010",
						 "100101100010000110101100",
						 "100101100010000011010110",
						 "100101100010000000000000",
						 "100101100001111100101010",
						 "100101100010101110110100",
						 "100101100010101011011110",
						 "100101100010101000001000",
						 "100101100010100100110010",
						 "100101100010100001011100",
						 "100101100010011110000110",
						 "100101100010011010110000",
						 "100101100010010111011010",
						 "100101100010010100000100",
						 "100101100010010000101110",
						 "100101100010001101011000",
						 "100101100010001010000010",
						 "100101100010000110101100",
						 "100101100010000011010110",
						 "100101100010000000000000",
						 "100101100001111100101010",
						 "100101100000001011110110",
						 "100101100000001000100000",
						 "100101100000000101001010",
						 "100101100000000001110100",
						 "100101011111111110011110",
						 "100101011111111011001000",
						 "100101011111110111110010",
						 "100101011111110100011100",
						 "100101011111110001000110",
						 "100101011111101101110000",
						 "100101011111101010011010",
						 "100101011111100111000100",
						 "100101011111100011101110",
						 "100101011111100000011000",
						 "100101011111011101000010",
						 "100101011111011001101100",
						 "100101100000001011110110",
						 "100101100000001000100000",
						 "100101100000000101001010",
						 "100101100000000001110100",
						 "100101011111111110011110",
						 "100101011111111011001000",
						 "100101011111110111110010",
						 "100101011111110100011100",
						 "100101011111110001000110",
						 "100101011111101101110000",
						 "100101011111101010011010",
						 "100101011111100111000100",
						 "100101011111100011101110",
						 "100101011111100000011000",
						 "100101011111011101000010",
						 "100101011111011001101100",
						 "100101100000001011110110",
						 "100101100000001000100000",
						 "100101100000000101001010",
						 "100101100000000001110100",
						 "100101011111111110011110",
						 "100101011111111011001000",
						 "100101011111110111110010",
						 "100101011111110100011100",
						 "100101011111110001000110",
						 "100101011111101101110000",
						 "100101011111101010011010",
						 "100101011111100111000100",
						 "100101011111100011101110",
						 "100101011111100000011000",
						 "100101011111011101000010",
						 "100101011111011001101100",
						 "100101011101101001000111",
						 "100101011101100101110000",
						 "100101011101100010011001",
						 "100101011101011111000010",
						 "100101011101011011101011",
						 "100101011101011000010100",
						 "100101011101010100111101",
						 "100101011101010001100110",
						 "100101011101001110001111",
						 "100101011101001010111000",
						 "100101011101000111100001",
						 "100101011101000100001010",
						 "100101011101000000110011",
						 "100101011100111101011100",
						 "100101011100111010000101",
						 "100101011100110110101110",
						 "100101011101101001000111",
						 "100101011101100101110000",
						 "100101011101100010011001",
						 "100101011101011111000010",
						 "100101011101011011101011",
						 "100101011101011000010100",
						 "100101011101010100111101",
						 "100101011101010001100110",
						 "100101011101001110001111",
						 "100101011101001010111000",
						 "100101011101000111100001",
						 "100101011101000100001010",
						 "100101011101000000110011",
						 "100101011100111101011100",
						 "100101011100111010000101",
						 "100101011100110110101110",
						 "100101011101101001000111",
						 "100101011101100101110000",
						 "100101011101100010011001",
						 "100101011101011111000010",
						 "100101011101011011101011",
						 "100101011101011000010100",
						 "100101011101010100111101",
						 "100101011101010001100110",
						 "100101011101001110001111",
						 "100101011101001010111000",
						 "100101011101000111100001",
						 "100101011101000100001010",
						 "100101011101000000110011",
						 "100101011100111101011100",
						 "100101011100111010000101",
						 "100101011100110110101110",
						 "100101011011000110001001",
						 "100101011011000010110010",
						 "100101011010111111011011",
						 "100101011010111100000100",
						 "100101011010111000101101",
						 "100101011010110101010110",
						 "100101011010110001111111",
						 "100101011010101110101000",
						 "100101011010101011010001",
						 "100101011010100111111010",
						 "100101011010100100100011",
						 "100101011010100001001100",
						 "100101011010011101110101",
						 "100101011010011010011110",
						 "100101011010010111000111",
						 "100101011010010011110000",
						 "100101011011000110011000",
						 "100101011011000011000000",
						 "100101011010111111101000",
						 "100101011010111100010000",
						 "100101011010111000111000",
						 "100101011010110101100000",
						 "100101011010110010001000",
						 "100101011010101110110000",
						 "100101011010101011011000",
						 "100101011010101000000000",
						 "100101011010100100101000",
						 "100101011010100001010000",
						 "100101011010011101111000",
						 "100101011010011010100000",
						 "100101011010010111001000",
						 "100101011010010011110000",
						 "100101011011000110011000",
						 "100101011011000011000000",
						 "100101011010111111101000",
						 "100101011010111100010000",
						 "100101011010111000111000",
						 "100101011010110101100000",
						 "100101011010110010001000",
						 "100101011010101110110000",
						 "100101011010101011011000",
						 "100101011010101000000000",
						 "100101011010100100101000",
						 "100101011010100001010000",
						 "100101011010011101111000",
						 "100101011010011010100000",
						 "100101011010010111001000",
						 "100101011010010011110000",
						 "100101011000100011011010",
						 "100101011000100000000010",
						 "100101011000011100101010",
						 "100101011000011001010010",
						 "100101011000010101111010",
						 "100101011000010010100010",
						 "100101011000001111001010",
						 "100101011000001011110010",
						 "100101011000001000011010",
						 "100101011000000101000010",
						 "100101011000000001101010",
						 "100101010111111110010010",
						 "100101010111111010111010",
						 "100101010111110111100010",
						 "100101010111110100001010",
						 "100101010111110000110010",
						 "100101011000100011011010",
						 "100101011000100000000010",
						 "100101011000011100101010",
						 "100101011000011001010010",
						 "100101011000010101111010",
						 "100101011000010010100010",
						 "100101011000001111001010",
						 "100101011000001011110010",
						 "100101011000001000011010",
						 "100101011000000101000010",
						 "100101011000000001101010",
						 "100101010111111110010010",
						 "100101010111111010111010",
						 "100101010111110111100010",
						 "100101010111110100001010",
						 "100101010111110000110010",
						 "100101011000100011011010",
						 "100101011000100000000010",
						 "100101011000011100101010",
						 "100101011000011001010010",
						 "100101011000010101111010",
						 "100101011000010010100010",
						 "100101011000001111001010",
						 "100101011000001011110010",
						 "100101011000001000011010",
						 "100101011000000101000010",
						 "100101011000000001101010",
						 "100101010111111110010010",
						 "100101010111111010111010",
						 "100101010111110111100010",
						 "100101010111110100001010",
						 "100101010111110000110010",
						 "100101010110000000101011",
						 "100101010101111101010010",
						 "100101010101111001111001",
						 "100101010101110110100000",
						 "100101010101110011000111",
						 "100101010101101111101110",
						 "100101010101101100010101",
						 "100101010101101000111100",
						 "100101010101100101100011",
						 "100101010101100010001010",
						 "100101010101011110110001",
						 "100101010101011011011000",
						 "100101010101010111111111",
						 "100101010101010100100110",
						 "100101010101010001001101",
						 "100101010101001101110100",
						 "100101010110000000101011",
						 "100101010101111101010010",
						 "100101010101111001111001",
						 "100101010101110110100000",
						 "100101010101110011000111",
						 "100101010101101111101110",
						 "100101010101101100010101",
						 "100101010101101000111100",
						 "100101010101100101100011",
						 "100101010101100010001010",
						 "100101010101011110110001",
						 "100101010101011011011000",
						 "100101010101010111111111",
						 "100101010101010100100110",
						 "100101010101010001001101",
						 "100101010101001101110100",
						 "100101010110000000101011",
						 "100101010101111101010010",
						 "100101010101111001111001",
						 "100101010101110110100000",
						 "100101010101110011000111",
						 "100101010101101111101110",
						 "100101010101101100010101",
						 "100101010101101000111100",
						 "100101010101100101100011",
						 "100101010101100010001010",
						 "100101010101011110110001",
						 "100101010101011011011000",
						 "100101010101010111111111",
						 "100101010101010100100110",
						 "100101010101010001001101",
						 "100101010101001101110100",
						 "100101010011011101101101",
						 "100101010011011010010100",
						 "100101010011010110111011",
						 "100101010011010011100010",
						 "100101010011010000001001",
						 "100101010011001100110000",
						 "100101010011001001010111",
						 "100101010011000101111110",
						 "100101010011000010100101",
						 "100101010010111111001100",
						 "100101010010111011110011",
						 "100101010010111000011010",
						 "100101010010110101000001",
						 "100101010010110001101000",
						 "100101010010101110001111",
						 "100101010010101010110110",
						 "100101010011011101101101",
						 "100101010011011010010100",
						 "100101010011010110111011",
						 "100101010011010011100010",
						 "100101010011010000001001",
						 "100101010011001100110000",
						 "100101010011001001010111",
						 "100101010011000101111110",
						 "100101010011000010100101",
						 "100101010010111111001100",
						 "100101010010111011110011",
						 "100101010010111000011010",
						 "100101010010110101000001",
						 "100101010010110001101000",
						 "100101010010101110001111",
						 "100101010010101010110110",
						 "100101010011011101111100",
						 "100101010011011010100010",
						 "100101010011010111001000",
						 "100101010011010011101110",
						 "100101010011010000010100",
						 "100101010011001100111010",
						 "100101010011001001100000",
						 "100101010011000110000110",
						 "100101010011000010101100",
						 "100101010010111111010010",
						 "100101010010111011111000",
						 "100101010010111000011110",
						 "100101010010110101000100",
						 "100101010010110001101010",
						 "100101010010101110010000",
						 "100101010010101010110110",
						 "100101010000111010111110",
						 "100101010000110111100100",
						 "100101010000110100001010",
						 "100101010000110000110000",
						 "100101010000101101010110",
						 "100101010000101001111100",
						 "100101010000100110100010",
						 "100101010000100011001000",
						 "100101010000011111101110",
						 "100101010000011100010100",
						 "100101010000011000111010",
						 "100101010000010101100000",
						 "100101010000010010000110",
						 "100101010000001110101100",
						 "100101010000001011010010",
						 "100101010000000111111000",
						 "100101010000111010111110",
						 "100101010000110111100100",
						 "100101010000110100001010",
						 "100101010000110000110000",
						 "100101010000101101010110",
						 "100101010000101001111100",
						 "100101010000100110100010",
						 "100101010000100011001000",
						 "100101010000011111101110",
						 "100101010000011100010100",
						 "100101010000011000111010",
						 "100101010000010101100000",
						 "100101010000010010000110",
						 "100101010000001110101100",
						 "100101010000001011010010",
						 "100101010000000111111000",
						 "100101010000111010111110",
						 "100101010000110111100100",
						 "100101010000110100001010",
						 "100101010000110000110000",
						 "100101010000101101010110",
						 "100101010000101001111100",
						 "100101010000100110100010",
						 "100101010000100011001000",
						 "100101010000011111101110",
						 "100101010000011100010100",
						 "100101010000011000111010",
						 "100101010000010101100000",
						 "100101010000010010000110",
						 "100101010000001110101100",
						 "100101010000001011010010",
						 "100101010000000111111000",
						 "100101001110011000000000",
						 "100101001110010100100110",
						 "100101001110010001001100",
						 "100101001110001101110010",
						 "100101001110001010011000",
						 "100101001110000110111110",
						 "100101001110000011100100",
						 "100101001110000000001010",
						 "100101001101111100110000",
						 "100101001101111001010110",
						 "100101001101110101111100",
						 "100101001101110010100010",
						 "100101001101101111001000",
						 "100101001101101011101110",
						 "100101001101101000010100",
						 "100101001101100100111010",
						 "100101001110011000001111",
						 "100101001110010100110100",
						 "100101001110010001011001",
						 "100101001110001101111110",
						 "100101001110001010100011",
						 "100101001110000111001000",
						 "100101001110000011101101",
						 "100101001110000000010010",
						 "100101001101111100110111",
						 "100101001101111001011100",
						 "100101001101110110000001",
						 "100101001101110010100110",
						 "100101001101101111001011",
						 "100101001101101011110000",
						 "100101001101101000010101",
						 "100101001101100100111010",
						 "100101001110011000001111",
						 "100101001110010100110100",
						 "100101001110010001011001",
						 "100101001110001101111110",
						 "100101001110001010100011",
						 "100101001110000111001000",
						 "100101001110000011101101",
						 "100101001110000000010010",
						 "100101001101111100110111",
						 "100101001101111001011100",
						 "100101001101110110000001",
						 "100101001101110010100110",
						 "100101001101101111001011",
						 "100101001101101011110000",
						 "100101001101101000010101",
						 "100101001101100100111010",
						 "100101001011110101010001",
						 "100101001011110001110110",
						 "100101001011101110011011",
						 "100101001011101011000000",
						 "100101001011100111100101",
						 "100101001011100100001010",
						 "100101001011100000101111",
						 "100101001011011101010100",
						 "100101001011011001111001",
						 "100101001011010110011110",
						 "100101001011010011000011",
						 "100101001011001111101000",
						 "100101001011001100001101",
						 "100101001011001000110010",
						 "100101001011000101010111",
						 "100101001011000001111100",
						 "100101001011110101010001",
						 "100101001011110001110110",
						 "100101001011101110011011",
						 "100101001011101011000000",
						 "100101001011100111100101",
						 "100101001011100100001010",
						 "100101001011100000101111",
						 "100101001011011101010100",
						 "100101001011011001111001",
						 "100101001011010110011110",
						 "100101001011010011000011",
						 "100101001011001111101000",
						 "100101001011001100001101",
						 "100101001011001000110010",
						 "100101001011000101010111",
						 "100101001011000001111100",
						 "100101001011110101010001",
						 "100101001011110001110110",
						 "100101001011101110011011",
						 "100101001011101011000000",
						 "100101001011100111100101",
						 "100101001011100100001010",
						 "100101001011100000101111",
						 "100101001011011101010100",
						 "100101001011011001111001",
						 "100101001011010110011110",
						 "100101001011010011000011",
						 "100101001011001111101000",
						 "100101001011001100001101",
						 "100101001011001000110010",
						 "100101001011000101010111",
						 "100101001011000001111100",
						 "100101001001010010100010",
						 "100101001001001111000110",
						 "100101001001001011101010",
						 "100101001001001000001110",
						 "100101001001000100110010",
						 "100101001001000001010110",
						 "100101001000111101111010",
						 "100101001000111010011110",
						 "100101001000110111000010",
						 "100101001000110011100110",
						 "100101001000110000001010",
						 "100101001000101100101110",
						 "100101001000101001010010",
						 "100101001000100101110110",
						 "100101001000100010011010",
						 "100101001000011110111110",
						 "100101001001010010100010",
						 "100101001001001111000110",
						 "100101001001001011101010",
						 "100101001001001000001110",
						 "100101001001000100110010",
						 "100101001001000001010110",
						 "100101001000111101111010",
						 "100101001000111010011110",
						 "100101001000110111000010",
						 "100101001000110011100110",
						 "100101001000110000001010",
						 "100101001000101100101110",
						 "100101001000101001010010",
						 "100101001000100101110110",
						 "100101001000100010011010",
						 "100101001000011110111110",
						 "100101001001010010100010",
						 "100101001001001111000110",
						 "100101001001001011101010",
						 "100101001001001000001110",
						 "100101001001000100110010",
						 "100101001001000001010110",
						 "100101001000111101111010",
						 "100101001000111010011110",
						 "100101001000110111000010",
						 "100101001000110011100110",
						 "100101001000110000001010",
						 "100101001000101100101110",
						 "100101001000101001010010",
						 "100101001000100101110110",
						 "100101001000100010011010",
						 "100101001000011110111110",
						 "100101000110101111100100",
						 "100101000110101100001000",
						 "100101000110101000101100",
						 "100101000110100101010000",
						 "100101000110100001110100",
						 "100101000110011110011000",
						 "100101000110011010111100",
						 "100101000110010111100000",
						 "100101000110010100000100",
						 "100101000110010000101000",
						 "100101000110001101001100",
						 "100101000110001001110000",
						 "100101000110000110010100",
						 "100101000110000010111000",
						 "100101000101111111011100",
						 "100101000101111100000000",
						 "100101000110101111100100",
						 "100101000110101100001000",
						 "100101000110101000101100",
						 "100101000110100101010000",
						 "100101000110100001110100",
						 "100101000110011110011000",
						 "100101000110011010111100",
						 "100101000110010111100000",
						 "100101000110010100000100",
						 "100101000110010000101000",
						 "100101000110001101001100",
						 "100101000110001001110000",
						 "100101000110000110010100",
						 "100101000110000010111000",
						 "100101000101111111011100",
						 "100101000101111100000000",
						 "100101000110101111110011",
						 "100101000110101100010110",
						 "100101000110101000111001",
						 "100101000110100101011100",
						 "100101000110100001111111",
						 "100101000110011110100010",
						 "100101000110011011000101",
						 "100101000110010111101000",
						 "100101000110010100001011",
						 "100101000110010000101110",
						 "100101000110001101010001",
						 "100101000110001001110100",
						 "100101000110000110010111",
						 "100101000110000010111010",
						 "100101000101111111011101",
						 "100101000101111100000000",
						 "100101000100001100110101",
						 "100101000100001001011000",
						 "100101000100000101111011",
						 "100101000100000010011110",
						 "100101000011111111000001",
						 "100101000011111011100100",
						 "100101000011111000000111",
						 "100101000011110100101010",
						 "100101000011110001001101",
						 "100101000011101101110000",
						 "100101000011101010010011",
						 "100101000011100110110110",
						 "100101000011100011011001",
						 "100101000011011111111100",
						 "100101000011011100011111",
						 "100101000011011001000010",
						 "100101000100001100110101",
						 "100101000100001001011000",
						 "100101000100000101111011",
						 "100101000100000010011110",
						 "100101000011111111000001",
						 "100101000011111011100100",
						 "100101000011111000000111",
						 "100101000011110100101010",
						 "100101000011110001001101",
						 "100101000011101101110000",
						 "100101000011101010010011",
						 "100101000011100110110110",
						 "100101000011100011011001",
						 "100101000011011111111100",
						 "100101000011011100011111",
						 "100101000011011001000010",
						 "100101000100001100110101",
						 "100101000100001001011000",
						 "100101000100000101111011",
						 "100101000100000010011110",
						 "100101000011111111000001",
						 "100101000011111011100100",
						 "100101000011111000000111",
						 "100101000011110100101010",
						 "100101000011110001001101",
						 "100101000011101101110000",
						 "100101000011101010010011",
						 "100101000011100110110110",
						 "100101000011100011011001",
						 "100101000011011111111100",
						 "100101000011011100011111",
						 "100101000011011001000010",
						 "100101000001101001110111",
						 "100101000001100110011010",
						 "100101000001100010111101",
						 "100101000001011111100000",
						 "100101000001011100000011",
						 "100101000001011000100110",
						 "100101000001010101001001",
						 "100101000001010001101100",
						 "100101000001001110001111",
						 "100101000001001010110010",
						 "100101000001000111010101",
						 "100101000001000011111000",
						 "100101000001000000011011",
						 "100101000000111100111110",
						 "100101000000111001100001",
						 "100101000000110110000100",
						 "100101000001101010000110",
						 "100101000001100110101000",
						 "100101000001100011001010",
						 "100101000001011111101100",
						 "100101000001011100001110",
						 "100101000001011000110000",
						 "100101000001010101010010",
						 "100101000001010001110100",
						 "100101000001001110010110",
						 "100101000001001010111000",
						 "100101000001000111011010",
						 "100101000001000011111100",
						 "100101000001000000011110",
						 "100101000000111101000000",
						 "100101000000111001100010",
						 "100101000000110110000100",
						 "100101000001101010000110",
						 "100101000001100110101000",
						 "100101000001100011001010",
						 "100101000001011111101100",
						 "100101000001011100001110",
						 "100101000001011000110000",
						 "100101000001010101010010",
						 "100101000001010001110100",
						 "100101000001001110010110",
						 "100101000001001010111000",
						 "100101000001000111011010",
						 "100101000001000011111100",
						 "100101000001000000011110",
						 "100101000000111101000000",
						 "100101000000111001100010",
						 "100101000000110110000100",
						 "100100111111000111001000",
						 "100100111111000011101010",
						 "100100111111000000001100",
						 "100100111110111100101110",
						 "100100111110111001010000",
						 "100100111110110101110010",
						 "100100111110110010010100",
						 "100100111110101110110110",
						 "100100111110101011011000",
						 "100100111110100111111010",
						 "100100111110100100011100",
						 "100100111110100000111110",
						 "100100111110011101100000",
						 "100100111110011010000010",
						 "100100111110010110100100",
						 "100100111110010011000110",
						 "100100111111000111001000",
						 "100100111111000011101010",
						 "100100111111000000001100",
						 "100100111110111100101110",
						 "100100111110111001010000",
						 "100100111110110101110010",
						 "100100111110110010010100",
						 "100100111110101110110110",
						 "100100111110101011011000",
						 "100100111110100111111010",
						 "100100111110100100011100",
						 "100100111110100000111110",
						 "100100111110011101100000",
						 "100100111110011010000010",
						 "100100111110010110100100",
						 "100100111110010011000110",
						 "100100111111000111001000",
						 "100100111111000011101010",
						 "100100111111000000001100",
						 "100100111110111100101110",
						 "100100111110111001010000",
						 "100100111110110101110010",
						 "100100111110110010010100",
						 "100100111110101110110110",
						 "100100111110101011011000",
						 "100100111110100111111010",
						 "100100111110100100011100",
						 "100100111110100000111110",
						 "100100111110011101100000",
						 "100100111110011010000010",
						 "100100111110010110100100",
						 "100100111110010011000110",
						 "100100111100100100011001",
						 "100100111100100000111010",
						 "100100111100011101011011",
						 "100100111100011001111100",
						 "100100111100010110011101",
						 "100100111100010010111110",
						 "100100111100001111011111",
						 "100100111100001100000000",
						 "100100111100001000100001",
						 "100100111100000101000010",
						 "100100111100000001100011",
						 "100100111011111110000100",
						 "100100111011111010100101",
						 "100100111011110111000110",
						 "100100111011110011100111",
						 "100100111011110000001000",
						 "100100111100100100011001",
						 "100100111100100000111010",
						 "100100111100011101011011",
						 "100100111100011001111100",
						 "100100111100010110011101",
						 "100100111100010010111110",
						 "100100111100001111011111",
						 "100100111100001100000000",
						 "100100111100001000100001",
						 "100100111100000101000010",
						 "100100111100000001100011",
						 "100100111011111110000100",
						 "100100111011111010100101",
						 "100100111011110111000110",
						 "100100111011110011100111",
						 "100100111011110000001000",
						 "100100111100100100011001",
						 "100100111100100000111010",
						 "100100111100011101011011",
						 "100100111100011001111100",
						 "100100111100010110011101",
						 "100100111100010010111110",
						 "100100111100001111011111",
						 "100100111100001100000000",
						 "100100111100001000100001",
						 "100100111100000101000010",
						 "100100111100000001100011",
						 "100100111011111110000100",
						 "100100111011111010100101",
						 "100100111011110111000110",
						 "100100111011110011100111",
						 "100100111011110000001000",
						 "100100111010000001011011",
						 "100100111001111101111100",
						 "100100111001111010011101",
						 "100100111001110110111110",
						 "100100111001110011011111",
						 "100100111001110000000000",
						 "100100111001101100100001",
						 "100100111001101001000010",
						 "100100111001100101100011",
						 "100100111001100010000100",
						 "100100111001011110100101",
						 "100100111001011011000110",
						 "100100111001010111100111",
						 "100100111001010100001000",
						 "100100111001010000101001",
						 "100100111001001101001010",
						 "100100111010000001011011",
						 "100100111001111101111100",
						 "100100111001111010011101",
						 "100100111001110110111110",
						 "100100111001110011011111",
						 "100100111001110000000000",
						 "100100111001101100100001",
						 "100100111001101001000010",
						 "100100111001100101100011",
						 "100100111001100010000100",
						 "100100111001011110100101",
						 "100100111001011011000110",
						 "100100111001010111100111",
						 "100100111001010100001000",
						 "100100111001010000101001",
						 "100100111001001101001010",
						 "100100111010000001011011",
						 "100100111001111101111100",
						 "100100111001111010011101",
						 "100100111001110110111110",
						 "100100111001110011011111",
						 "100100111001110000000000",
						 "100100111001101100100001",
						 "100100111001101001000010",
						 "100100111001100101100011",
						 "100100111001100010000100",
						 "100100111001011110100101",
						 "100100111001011011000110",
						 "100100111001010111100111",
						 "100100111001010100001000",
						 "100100111001010000101001",
						 "100100111001001101001010",
						 "100100110111011110101100",
						 "100100110111011011001100",
						 "100100110111010111101100",
						 "100100110111010100001100",
						 "100100110111010000101100",
						 "100100110111001101001100",
						 "100100110111001001101100",
						 "100100110111000110001100",
						 "100100110111000010101100",
						 "100100110110111111001100",
						 "100100110110111011101100",
						 "100100110110111000001100",
						 "100100110110110100101100",
						 "100100110110110001001100",
						 "100100110110101101101100",
						 "100100110110101010001100",
						 "100100110111011110101100",
						 "100100110111011011001100",
						 "100100110111010111101100",
						 "100100110111010100001100",
						 "100100110111010000101100",
						 "100100110111001101001100",
						 "100100110111001001101100",
						 "100100110111000110001100",
						 "100100110111000010101100",
						 "100100110110111111001100",
						 "100100110110111011101100",
						 "100100110110111000001100",
						 "100100110110110100101100",
						 "100100110110110001001100",
						 "100100110110101101101100",
						 "100100110110101010001100",
						 "100100110111011110101100",
						 "100100110111011011001100",
						 "100100110111010111101100",
						 "100100110111010100001100",
						 "100100110111010000101100",
						 "100100110111001101001100",
						 "100100110111001001101100",
						 "100100110111000110001100",
						 "100100110111000010101100",
						 "100100110110111111001100",
						 "100100110110111011101100",
						 "100100110110111000001100",
						 "100100110110110100101100",
						 "100100110110110001001100",
						 "100100110110101101101100",
						 "100100110110101010001100",
						 "100100110100111011101110",
						 "100100110100111000001110",
						 "100100110100110100101110",
						 "100100110100110001001110",
						 "100100110100101101101110",
						 "100100110100101010001110",
						 "100100110100100110101110",
						 "100100110100100011001110",
						 "100100110100011111101110",
						 "100100110100011100001110",
						 "100100110100011000101110",
						 "100100110100010101001110",
						 "100100110100010001101110",
						 "100100110100001110001110",
						 "100100110100001010101110",
						 "100100110100000111001110",
						 "100100110100111011101110",
						 "100100110100111000001110",
						 "100100110100110100101110",
						 "100100110100110001001110",
						 "100100110100101101101110",
						 "100100110100101010001110",
						 "100100110100100110101110",
						 "100100110100100011001110",
						 "100100110100011111101110",
						 "100100110100011100001110",
						 "100100110100011000101110",
						 "100100110100010101001110",
						 "100100110100010001101110",
						 "100100110100001110001110",
						 "100100110100001010101110",
						 "100100110100000111001110",
						 "100100110100111011111101",
						 "100100110100111000011100",
						 "100100110100110100111011",
						 "100100110100110001011010",
						 "100100110100101101111001",
						 "100100110100101010011000",
						 "100100110100100110110111",
						 "100100110100100011010110",
						 "100100110100011111110101",
						 "100100110100011100010100",
						 "100100110100011000110011",
						 "100100110100010101010010",
						 "100100110100010001110001",
						 "100100110100001110010000",
						 "100100110100001010101111",
						 "100100110100000111001110",
						 "100100110010011000111111",
						 "100100110010010101011110",
						 "100100110010010001111101",
						 "100100110010001110011100",
						 "100100110010001010111011",
						 "100100110010000111011010",
						 "100100110010000011111001",
						 "100100110010000000011000",
						 "100100110001111100110111",
						 "100100110001111001010110",
						 "100100110001110101110101",
						 "100100110001110010010100",
						 "100100110001101110110011",
						 "100100110001101011010010",
						 "100100110001100111110001",
						 "100100110001100100010000",
						 "100100110010011000111111",
						 "100100110010010101011110",
						 "100100110010010001111101",
						 "100100110010001110011100",
						 "100100110010001010111011",
						 "100100110010000111011010",
						 "100100110010000011111001",
						 "100100110010000000011000",
						 "100100110001111100110111",
						 "100100110001111001010110",
						 "100100110001110101110101",
						 "100100110001110010010100",
						 "100100110001101110110011",
						 "100100110001101011010010",
						 "100100110001100111110001",
						 "100100110001100100010000",
						 "100100110010011000111111",
						 "100100110010010101011110",
						 "100100110010010001111101",
						 "100100110010001110011100",
						 "100100110010001010111011",
						 "100100110010000111011010",
						 "100100110010000011111001",
						 "100100110010000000011000",
						 "100100110001111100110111",
						 "100100110001111001010110",
						 "100100110001110101110101",
						 "100100110001110010010100",
						 "100100110001101110110011",
						 "100100110001101011010010",
						 "100100110001100111110001",
						 "100100110001100100010000",
						 "100100101111110110000001",
						 "100100101111110010100000",
						 "100100101111101110111111",
						 "100100101111101011011110",
						 "100100101111100111111101",
						 "100100101111100100011100",
						 "100100101111100000111011",
						 "100100101111011101011010",
						 "100100101111011001111001",
						 "100100101111010110011000",
						 "100100101111010010110111",
						 "100100101111001111010110",
						 "100100101111001011110101",
						 "100100101111001000010100",
						 "100100101111000100110011",
						 "100100101111000001010010",
						 "100100101111110110010000",
						 "100100101111110010101110",
						 "100100101111101111001100",
						 "100100101111101011101010",
						 "100100101111101000001000",
						 "100100101111100100100110",
						 "100100101111100001000100",
						 "100100101111011101100010",
						 "100100101111011010000000",
						 "100100101111010110011110",
						 "100100101111010010111100",
						 "100100101111001111011010",
						 "100100101111001011111000",
						 "100100101111001000010110",
						 "100100101111000100110100",
						 "100100101111000001010010",
						 "100100101101010011010010",
						 "100100101101001111110000",
						 "100100101101001100001110",
						 "100100101101001000101100",
						 "100100101101000101001010",
						 "100100101101000001101000",
						 "100100101100111110000110",
						 "100100101100111010100100",
						 "100100101100110111000010",
						 "100100101100110011100000",
						 "100100101100101111111110",
						 "100100101100101100011100",
						 "100100101100101000111010",
						 "100100101100100101011000",
						 "100100101100100001110110",
						 "100100101100011110010100",
						 "100100101101010011010010",
						 "100100101101001111110000",
						 "100100101101001100001110",
						 "100100101101001000101100",
						 "100100101101000101001010",
						 "100100101101000001101000",
						 "100100101100111110000110",
						 "100100101100111010100100",
						 "100100101100110111000010",
						 "100100101100110011100000",
						 "100100101100101111111110",
						 "100100101100101100011100",
						 "100100101100101000111010",
						 "100100101100100101011000",
						 "100100101100100001110110",
						 "100100101100011110010100",
						 "100100101101010011010010",
						 "100100101101001111110000",
						 "100100101101001100001110",
						 "100100101101001000101100",
						 "100100101101000101001010",
						 "100100101101000001101000",
						 "100100101100111110000110",
						 "100100101100111010100100",
						 "100100101100110111000010",
						 "100100101100110011100000",
						 "100100101100101111111110",
						 "100100101100101100011100",
						 "100100101100101000111010",
						 "100100101100100101011000",
						 "100100101100100001110110",
						 "100100101100011110010100",
						 "100100101010110000010100",
						 "100100101010101100110010",
						 "100100101010101001010000",
						 "100100101010100101101110",
						 "100100101010100010001100",
						 "100100101010011110101010",
						 "100100101010011011001000",
						 "100100101010010111100110",
						 "100100101010010100000100",
						 "100100101010010000100010",
						 "100100101010001101000000",
						 "100100101010001001011110",
						 "100100101010000101111100",
						 "100100101010000010011010",
						 "100100101001111110111000",
						 "100100101001111011010110",
						 "100100101010110000010100",
						 "100100101010101100110010",
						 "100100101010101001010000",
						 "100100101010100101101110",
						 "100100101010100010001100",
						 "100100101010011110101010",
						 "100100101010011011001000",
						 "100100101010010111100110",
						 "100100101010010100000100",
						 "100100101010010000100010",
						 "100100101010001101000000",
						 "100100101010001001011110",
						 "100100101010000101111100",
						 "100100101010000010011010",
						 "100100101001111110111000",
						 "100100101001111011010110",
						 "100100101010110000100011",
						 "100100101010101101000000",
						 "100100101010101001011101",
						 "100100101010100101111010",
						 "100100101010100010010111",
						 "100100101010011110110100",
						 "100100101010011011010001",
						 "100100101010010111101110",
						 "100100101010010100001011",
						 "100100101010010000101000",
						 "100100101010001101000101",
						 "100100101010001001100010",
						 "100100101010000101111111",
						 "100100101010000010011100",
						 "100100101001111110111001",
						 "100100101001111011010110",
						 "100100101000001101100101",
						 "100100101000001010000010",
						 "100100101000000110011111",
						 "100100101000000010111100",
						 "100100100111111111011001",
						 "100100100111111011110110",
						 "100100100111111000010011",
						 "100100100111110100110000",
						 "100100100111110001001101",
						 "100100100111101101101010",
						 "100100100111101010000111",
						 "100100100111100110100100",
						 "100100100111100011000001",
						 "100100100111011111011110",
						 "100100100111011011111011",
						 "100100100111011000011000",
						 "100100101000001101100101",
						 "100100101000001010000010",
						 "100100101000000110011111",
						 "100100101000000010111100",
						 "100100100111111111011001",
						 "100100100111111011110110",
						 "100100100111111000010011",
						 "100100100111110100110000",
						 "100100100111110001001101",
						 "100100100111101101101010",
						 "100100100111101010000111",
						 "100100100111100110100100",
						 "100100100111100011000001",
						 "100100100111011111011110",
						 "100100100111011011111011",
						 "100100100111011000011000",
						 "100100101000001101100101",
						 "100100101000001010000010",
						 "100100101000000110011111",
						 "100100101000000010111100",
						 "100100100111111111011001",
						 "100100100111111011110110",
						 "100100100111111000010011",
						 "100100100111110100110000",
						 "100100100111110001001101",
						 "100100100111101101101010",
						 "100100100111101010000111",
						 "100100100111100110100100",
						 "100100100111100011000001",
						 "100100100111011111011110",
						 "100100100111011011111011",
						 "100100100111011000011000",
						 "100100100101101010100111",
						 "100100100101100111000100",
						 "100100100101100011100001",
						 "100100100101011111111110",
						 "100100100101011100011011",
						 "100100100101011000111000",
						 "100100100101010101010101",
						 "100100100101010001110010",
						 "100100100101001110001111",
						 "100100100101001010101100",
						 "100100100101000111001001",
						 "100100100101000011100110",
						 "100100100101000000000011",
						 "100100100100111100100000",
						 "100100100100111000111101",
						 "100100100100110101011010",
						 "100100100101101010110110",
						 "100100100101100111010010",
						 "100100100101100011101110",
						 "100100100101100000001010",
						 "100100100101011100100110",
						 "100100100101011001000010",
						 "100100100101010101011110",
						 "100100100101010001111010",
						 "100100100101001110010110",
						 "100100100101001010110010",
						 "100100100101000111001110",
						 "100100100101000011101010",
						 "100100100101000000000110",
						 "100100100100111100100010",
						 "100100100100111000111110",
						 "100100100100110101011010",
						 "100100100101101010110110",
						 "100100100101100111010010",
						 "100100100101100011101110",
						 "100100100101100000001010",
						 "100100100101011100100110",
						 "100100100101011001000010",
						 "100100100101010101011110",
						 "100100100101010001111010",
						 "100100100101001110010110",
						 "100100100101001010110010",
						 "100100100101000111001110",
						 "100100100101000011101010",
						 "100100100101000000000110",
						 "100100100100111100100010",
						 "100100100100111000111110",
						 "100100100100110101011010",
						 "100100100011000111111000",
						 "100100100011000100010100",
						 "100100100011000000110000",
						 "100100100010111101001100",
						 "100100100010111001101000",
						 "100100100010110110000100",
						 "100100100010110010100000",
						 "100100100010101110111100",
						 "100100100010101011011000",
						 "100100100010100111110100",
						 "100100100010100100010000",
						 "100100100010100000101100",
						 "100100100010011101001000",
						 "100100100010011001100100",
						 "100100100010010110000000",
						 "100100100010010010011100",
						 "100100100011000111111000",
						 "100100100011000100010100",
						 "100100100011000000110000",
						 "100100100010111101001100",
						 "100100100010111001101000",
						 "100100100010110110000100",
						 "100100100010110010100000",
						 "100100100010101110111100",
						 "100100100010101011011000",
						 "100100100010100111110100",
						 "100100100010100100010000",
						 "100100100010100000101100",
						 "100100100010011101001000",
						 "100100100010011001100100",
						 "100100100010010110000000",
						 "100100100010010010011100",
						 "100100100011000111111000",
						 "100100100011000100010100",
						 "100100100011000000110000",
						 "100100100010111101001100",
						 "100100100010111001101000",
						 "100100100010110110000100",
						 "100100100010110010100000",
						 "100100100010101110111100",
						 "100100100010101011011000",
						 "100100100010100111110100",
						 "100100100010100100010000",
						 "100100100010100000101100",
						 "100100100010011101001000",
						 "100100100010011001100100",
						 "100100100010010110000000",
						 "100100100010010010011100",
						 "100100100000100100111010",
						 "100100100000100001010110",
						 "100100100000011101110010",
						 "100100100000011010001110",
						 "100100100000010110101010",
						 "100100100000010011000110",
						 "100100100000001111100010",
						 "100100100000001011111110",
						 "100100100000001000011010",
						 "100100100000000100110110",
						 "100100100000000001010010",
						 "100100011111111101101110",
						 "100100011111111010001010",
						 "100100011111110110100110",
						 "100100011111110011000010",
						 "100100011111101111011110",
						 "100100100000100101001001",
						 "100100100000100001100100",
						 "100100100000011101111111",
						 "100100100000011010011010",
						 "100100100000010110110101",
						 "100100100000010011010000",
						 "100100100000001111101011",
						 "100100100000001100000110",
						 "100100100000001000100001",
						 "100100100000000100111100",
						 "100100100000000001010111",
						 "100100011111111101110010",
						 "100100011111111010001101",
						 "100100011111110110101000",
						 "100100011111110011000011",
						 "100100011111101111011110",
						 "100100100000100101001001",
						 "100100100000100001100100",
						 "100100100000011101111111",
						 "100100100000011010011010",
						 "100100100000010110110101",
						 "100100100000010011010000",
						 "100100100000001111101011",
						 "100100100000001100000110",
						 "100100100000001000100001",
						 "100100100000000100111100",
						 "100100100000000001010111",
						 "100100011111111101110010",
						 "100100011111111010001101",
						 "100100011111110110101000",
						 "100100011111110011000011",
						 "100100011111101111011110",
						 "100100011110000010001011",
						 "100100011101111110100110",
						 "100100011101111011000001",
						 "100100011101110111011100",
						 "100100011101110011110111",
						 "100100011101110000010010",
						 "100100011101101100101101",
						 "100100011101101001001000",
						 "100100011101100101100011",
						 "100100011101100001111110",
						 "100100011101011110011001",
						 "100100011101011010110100",
						 "100100011101010111001111",
						 "100100011101010011101010",
						 "100100011101010000000101",
						 "100100011101001100100000",
						 "100100011110000010001011",
						 "100100011101111110100110",
						 "100100011101111011000001",
						 "100100011101110111011100",
						 "100100011101110011110111",
						 "100100011101110000010010",
						 "100100011101101100101101",
						 "100100011101101001001000",
						 "100100011101100101100011",
						 "100100011101100001111110",
						 "100100011101011110011001",
						 "100100011101011010110100",
						 "100100011101010111001111",
						 "100100011101010011101010",
						 "100100011101010000000101",
						 "100100011101001100100000",
						 "100100011011011111001101",
						 "100100011011011011101000",
						 "100100011011011000000011",
						 "100100011011010100011110",
						 "100100011011010000111001",
						 "100100011011001101010100",
						 "100100011011001001101111",
						 "100100011011000110001010",
						 "100100011011000010100101",
						 "100100011010111111000000",
						 "100100011010111011011011",
						 "100100011010110111110110",
						 "100100011010110100010001",
						 "100100011010110000101100",
						 "100100011010101101000111",
						 "100100011010101001100010",
						 "100100011011011111001101",
						 "100100011011011011101000",
						 "100100011011011000000011",
						 "100100011011010100011110",
						 "100100011011010000111001",
						 "100100011011001101010100",
						 "100100011011001001101111",
						 "100100011011000110001010",
						 "100100011011000010100101",
						 "100100011010111111000000",
						 "100100011010111011011011",
						 "100100011010110111110110",
						 "100100011010110100010001",
						 "100100011010110000101100",
						 "100100011010101101000111",
						 "100100011010101001100010",
						 "100100011011011111011100",
						 "100100011011011011110110",
						 "100100011011011000010000",
						 "100100011011010100101010",
						 "100100011011010001000100",
						 "100100011011001101011110",
						 "100100011011001001111000",
						 "100100011011000110010010",
						 "100100011011000010101100",
						 "100100011010111111000110",
						 "100100011010111011100000",
						 "100100011010110111111010",
						 "100100011010110100010100",
						 "100100011010110000101110",
						 "100100011010101101001000",
						 "100100011010101001100010",
						 "100100011000111100011110",
						 "100100011000111000111000",
						 "100100011000110101010010",
						 "100100011000110001101100",
						 "100100011000101110000110",
						 "100100011000101010100000",
						 "100100011000100110111010",
						 "100100011000100011010100",
						 "100100011000011111101110",
						 "100100011000011100001000",
						 "100100011000011000100010",
						 "100100011000010100111100",
						 "100100011000010001010110",
						 "100100011000001101110000",
						 "100100011000001010001010",
						 "100100011000000110100100",
						 "100100011000111100011110",
						 "100100011000111000111000",
						 "100100011000110101010010",
						 "100100011000110001101100",
						 "100100011000101110000110",
						 "100100011000101010100000",
						 "100100011000100110111010",
						 "100100011000100011010100",
						 "100100011000011111101110",
						 "100100011000011100001000",
						 "100100011000011000100010",
						 "100100011000010100111100",
						 "100100011000010001010110",
						 "100100011000001101110000",
						 "100100011000001010001010",
						 "100100011000000110100100",
						 "100100011000111100011110",
						 "100100011000111000111000",
						 "100100011000110101010010",
						 "100100011000110001101100",
						 "100100011000101110000110",
						 "100100011000101010100000",
						 "100100011000100110111010",
						 "100100011000100011010100",
						 "100100011000011111101110",
						 "100100011000011100001000",
						 "100100011000011000100010",
						 "100100011000010100111100",
						 "100100011000010001010110",
						 "100100011000001101110000",
						 "100100011000001010001010",
						 "100100011000000110100100",
						 "100100010110011001100000",
						 "100100010110010101111010",
						 "100100010110010010010100",
						 "100100010110001110101110",
						 "100100010110001011001000",
						 "100100010110000111100010",
						 "100100010110000011111100",
						 "100100010110000000010110",
						 "100100010101111100110000",
						 "100100010101111001001010",
						 "100100010101110101100100",
						 "100100010101110001111110",
						 "100100010101101110011000",
						 "100100010101101010110010",
						 "100100010101100111001100",
						 "100100010101100011100110",
						 "100100010110011001100000",
						 "100100010110010101111010",
						 "100100010110010010010100",
						 "100100010110001110101110",
						 "100100010110001011001000",
						 "100100010110000111100010",
						 "100100010110000011111100",
						 "100100010110000000010110",
						 "100100010101111100110000",
						 "100100010101111001001010",
						 "100100010101110101100100",
						 "100100010101110001111110",
						 "100100010101101110011000",
						 "100100010101101010110010",
						 "100100010101100111001100",
						 "100100010101100011100110",
						 "100100010110011001101111",
						 "100100010110010110001000",
						 "100100010110010010100001",
						 "100100010110001110111010",
						 "100100010110001011010011",
						 "100100010110000111101100",
						 "100100010110000100000101",
						 "100100010110000000011110",
						 "100100010101111100110111",
						 "100100010101111001010000",
						 "100100010101110101101001",
						 "100100010101110010000010",
						 "100100010101101110011011",
						 "100100010101101010110100",
						 "100100010101100111001101",
						 "100100010101100011100110",
						 "100100010011110110110001",
						 "100100010011110011001010",
						 "100100010011101111100011",
						 "100100010011101011111100",
						 "100100010011101000010101",
						 "100100010011100100101110",
						 "100100010011100001000111",
						 "100100010011011101100000",
						 "100100010011011001111001",
						 "100100010011010110010010",
						 "100100010011010010101011",
						 "100100010011001111000100",
						 "100100010011001011011101",
						 "100100010011000111110110",
						 "100100010011000100001111",
						 "100100010011000000101000",
						 "100100010011110110110001",
						 "100100010011110011001010",
						 "100100010011101111100011",
						 "100100010011101011111100",
						 "100100010011101000010101",
						 "100100010011100100101110",
						 "100100010011100001000111",
						 "100100010011011101100000",
						 "100100010011011001111001",
						 "100100010011010110010010",
						 "100100010011010010101011",
						 "100100010011001111000100",
						 "100100010011001011011101",
						 "100100010011000111110110",
						 "100100010011000100001111",
						 "100100010011000000101000",
						 "100100010011110110110001",
						 "100100010011110011001010",
						 "100100010011101111100011",
						 "100100010011101011111100",
						 "100100010011101000010101",
						 "100100010011100100101110",
						 "100100010011100001000111",
						 "100100010011011101100000",
						 "100100010011011001111001",
						 "100100010011010110010010",
						 "100100010011010010101011",
						 "100100010011001111000100",
						 "100100010011001011011101",
						 "100100010011000111110110",
						 "100100010011000100001111",
						 "100100010011000000101000",
						 "100100010001010011110011",
						 "100100010001010000001100",
						 "100100010001001100100101",
						 "100100010001001000111110",
						 "100100010001000101010111",
						 "100100010001000001110000",
						 "100100010000111110001001",
						 "100100010000111010100010",
						 "100100010000110110111011",
						 "100100010000110011010100",
						 "100100010000101111101101",
						 "100100010000101100000110",
						 "100100010000101000011111",
						 "100100010000100100111000",
						 "100100010000100001010001",
						 "100100010000011101101010",
						 "100100010001010011110011",
						 "100100010001010000001100",
						 "100100010001001100100101",
						 "100100010001001000111110",
						 "100100010001000101010111",
						 "100100010001000001110000",
						 "100100010000111110001001",
						 "100100010000111010100010",
						 "100100010000110110111011",
						 "100100010000110011010100",
						 "100100010000101111101101",
						 "100100010000101100000110",
						 "100100010000101000011111",
						 "100100010000100100111000",
						 "100100010000100001010001",
						 "100100010000011101101010",
						 "100100010001010100000010",
						 "100100010001010000011010",
						 "100100010001001100110010",
						 "100100010001001001001010",
						 "100100010001000101100010",
						 "100100010001000001111010",
						 "100100010000111110010010",
						 "100100010000111010101010",
						 "100100010000110111000010",
						 "100100010000110011011010",
						 "100100010000101111110010",
						 "100100010000101100001010",
						 "100100010000101000100010",
						 "100100010000100100111010",
						 "100100010000100001010010",
						 "100100010000011101101010",
						 "100100001110110001000100",
						 "100100001110101101011100",
						 "100100001110101001110100",
						 "100100001110100110001100",
						 "100100001110100010100100",
						 "100100001110011110111100",
						 "100100001110011011010100",
						 "100100001110010111101100",
						 "100100001110010100000100",
						 "100100001110010000011100",
						 "100100001110001100110100",
						 "100100001110001001001100",
						 "100100001110000101100100",
						 "100100001110000001111100",
						 "100100001101111110010100",
						 "100100001101111010101100",
						 "100100001110110001000100",
						 "100100001110101101011100",
						 "100100001110101001110100",
						 "100100001110100110001100",
						 "100100001110100010100100",
						 "100100001110011110111100",
						 "100100001110011011010100",
						 "100100001110010111101100",
						 "100100001110010100000100",
						 "100100001110010000011100",
						 "100100001110001100110100",
						 "100100001110001001001100",
						 "100100001110000101100100",
						 "100100001110000001111100",
						 "100100001101111110010100",
						 "100100001101111010101100",
						 "100100001100001110000110",
						 "100100001100001010011110",
						 "100100001100000110110110",
						 "100100001100000011001110",
						 "100100001011111111100110",
						 "100100001011111011111110",
						 "100100001011111000010110",
						 "100100001011110100101110",
						 "100100001011110001000110",
						 "100100001011101101011110",
						 "100100001011101001110110",
						 "100100001011100110001110",
						 "100100001011100010100110",
						 "100100001011011110111110",
						 "100100001011011011010110",
						 "100100001011010111101110",
						 "100100001100001110000110",
						 "100100001100001010011110",
						 "100100001100000110110110",
						 "100100001100000011001110",
						 "100100001011111111100110",
						 "100100001011111011111110",
						 "100100001011111000010110",
						 "100100001011110100101110",
						 "100100001011110001000110",
						 "100100001011101101011110",
						 "100100001011101001110110",
						 "100100001011100110001110",
						 "100100001011100010100110",
						 "100100001011011110111110",
						 "100100001011011011010110",
						 "100100001011010111101110",
						 "100100001100001110000110",
						 "100100001100001010011110",
						 "100100001100000110110110",
						 "100100001100000011001110",
						 "100100001011111111100110",
						 "100100001011111011111110",
						 "100100001011111000010110",
						 "100100001011110100101110",
						 "100100001011110001000110",
						 "100100001011101101011110",
						 "100100001011101001110110",
						 "100100001011100110001110",
						 "100100001011100010100110",
						 "100100001011011110111110",
						 "100100001011011011010110",
						 "100100001011010111101110",
						 "100100001001101011010111",
						 "100100001001100111101110",
						 "100100001001100100000101",
						 "100100001001100000011100",
						 "100100001001011100110011",
						 "100100001001011001001010",
						 "100100001001010101100001",
						 "100100001001010001111000",
						 "100100001001001110001111",
						 "100100001001001010100110",
						 "100100001001000110111101",
						 "100100001001000011010100",
						 "100100001000111111101011",
						 "100100001000111100000010",
						 "100100001000111000011001",
						 "100100001000110100110000",
						 "100100001001101011010111",
						 "100100001001100111101110",
						 "100100001001100100000101",
						 "100100001001100000011100",
						 "100100001001011100110011",
						 "100100001001011001001010",
						 "100100001001010101100001",
						 "100100001001010001111000",
						 "100100001001001110001111",
						 "100100001001001010100110",
						 "100100001001000110111101",
						 "100100001001000011010100",
						 "100100001000111111101011",
						 "100100001000111100000010",
						 "100100001000111000011001",
						 "100100001000110100110000",
						 "100100001001101011010111",
						 "100100001001100111101110",
						 "100100001001100100000101",
						 "100100001001100000011100",
						 "100100001001011100110011",
						 "100100001001011001001010",
						 "100100001001010101100001",
						 "100100001001010001111000",
						 "100100001001001110001111",
						 "100100001001001010100110",
						 "100100001001000110111101",
						 "100100001001000011010100",
						 "100100001000111111101011",
						 "100100001000111100000010",
						 "100100001000111000011001",
						 "100100001000110100110000",
						 "100100000111001000011001",
						 "100100000111000100110000",
						 "100100000111000001000111",
						 "100100000110111101011110",
						 "100100000110111001110101",
						 "100100000110110110001100",
						 "100100000110110010100011",
						 "100100000110101110111010",
						 "100100000110101011010001",
						 "100100000110100111101000",
						 "100100000110100011111111",
						 "100100000110100000010110",
						 "100100000110011100101101",
						 "100100000110011001000100",
						 "100100000110010101011011",
						 "100100000110010001110010",
						 "100100000111001000011001",
						 "100100000111000100110000",
						 "100100000111000001000111",
						 "100100000110111101011110",
						 "100100000110111001110101",
						 "100100000110110110001100",
						 "100100000110110010100011",
						 "100100000110101110111010",
						 "100100000110101011010001",
						 "100100000110100111101000",
						 "100100000110100011111111",
						 "100100000110100000010110",
						 "100100000110011100101101",
						 "100100000110011001000100",
						 "100100000110010101011011",
						 "100100000110010001110010",
						 "100100000111001000011001",
						 "100100000111000100110000",
						 "100100000111000001000111",
						 "100100000110111101011110",
						 "100100000110111001110101",
						 "100100000110110110001100",
						 "100100000110110010100011",
						 "100100000110101110111010",
						 "100100000110101011010001",
						 "100100000110100111101000",
						 "100100000110100011111111",
						 "100100000110100000010110",
						 "100100000110011100101101",
						 "100100000110011001000100",
						 "100100000110010101011011",
						 "100100000110010001110010",
						 "100100000100100101101010",
						 "100100000100100010000000",
						 "100100000100011110010110",
						 "100100000100011010101100",
						 "100100000100010111000010",
						 "100100000100010011011000",
						 "100100000100001111101110",
						 "100100000100001100000100",
						 "100100000100001000011010",
						 "100100000100000100110000",
						 "100100000100000001000110",
						 "100100000011111101011100",
						 "100100000011111001110010",
						 "100100000011110110001000",
						 "100100000011110010011110",
						 "100100000011101110110100",
						 "100100000100100101101010",
						 "100100000100100010000000",
						 "100100000100011110010110",
						 "100100000100011010101100",
						 "100100000100010111000010",
						 "100100000100010011011000",
						 "100100000100001111101110",
						 "100100000100001100000100",
						 "100100000100001000011010",
						 "100100000100000100110000",
						 "100100000100000001000110",
						 "100100000011111101011100",
						 "100100000011111001110010",
						 "100100000011110110001000",
						 "100100000011110010011110",
						 "100100000011101110110100",
						 "100100000100100101101010",
						 "100100000100100010000000",
						 "100100000100011110010110",
						 "100100000100011010101100",
						 "100100000100010111000010",
						 "100100000100010011011000",
						 "100100000100001111101110",
						 "100100000100001100000100",
						 "100100000100001000011010",
						 "100100000100000100110000",
						 "100100000100000001000110",
						 "100100000011111101011100",
						 "100100000011111001110010",
						 "100100000011110110001000",
						 "100100000011110010011110",
						 "100100000011101110110100",
						 "100100000010000010101100",
						 "100100000001111111000010",
						 "100100000001111011011000",
						 "100100000001110111101110",
						 "100100000001110100000100",
						 "100100000001110000011010",
						 "100100000001101100110000",
						 "100100000001101001000110",
						 "100100000001100101011100",
						 "100100000001100001110010",
						 "100100000001011110001000",
						 "100100000001011010011110",
						 "100100000001010110110100",
						 "100100000001010011001010",
						 "100100000001001111100000",
						 "100100000001001011110110",
						 "100100000010000010101100",
						 "100100000001111111000010",
						 "100100000001111011011000",
						 "100100000001110111101110",
						 "100100000001110100000100",
						 "100100000001110000011010",
						 "100100000001101100110000",
						 "100100000001101001000110",
						 "100100000001100101011100",
						 "100100000001100001110010",
						 "100100000001011110001000",
						 "100100000001011010011110",
						 "100100000001010110110100",
						 "100100000001010011001010",
						 "100100000001001111100000",
						 "100100000001001011110110",
						 "100011111111011111101110",
						 "100011111111011100000100",
						 "100011111111011000011010",
						 "100011111111010100110000",
						 "100011111111010001000110",
						 "100011111111001101011100",
						 "100011111111001001110010",
						 "100011111111000110001000",
						 "100011111111000010011110",
						 "100011111110111110110100",
						 "100011111110111011001010",
						 "100011111110110111100000",
						 "100011111110110011110110",
						 "100011111110110000001100",
						 "100011111110101100100010",
						 "100011111110101000111000",
						 "100011111111011111101110",
						 "100011111111011100000100",
						 "100011111111011000011010",
						 "100011111111010100110000",
						 "100011111111010001000110",
						 "100011111111001101011100",
						 "100011111111001001110010",
						 "100011111111000110001000",
						 "100011111111000010011110",
						 "100011111110111110110100",
						 "100011111110111011001010",
						 "100011111110110111100000",
						 "100011111110110011110110",
						 "100011111110110000001100",
						 "100011111110101100100010",
						 "100011111110101000111000",
						 "100011111111011111111101",
						 "100011111111011100010010",
						 "100011111111011000100111",
						 "100011111111010100111100",
						 "100011111111010001010001",
						 "100011111111001101100110",
						 "100011111111001001111011",
						 "100011111111000110010000",
						 "100011111111000010100101",
						 "100011111110111110111010",
						 "100011111110111011001111",
						 "100011111110110111100100",
						 "100011111110110011111001",
						 "100011111110110000001110",
						 "100011111110101100100011",
						 "100011111110101000111000",
						 "100011111100111100111111",
						 "100011111100111001010100",
						 "100011111100110101101001",
						 "100011111100110001111110",
						 "100011111100101110010011",
						 "100011111100101010101000",
						 "100011111100100110111101",
						 "100011111100100011010010",
						 "100011111100011111100111",
						 "100011111100011011111100",
						 "100011111100011000010001",
						 "100011111100010100100110",
						 "100011111100010000111011",
						 "100011111100001101010000",
						 "100011111100001001100101",
						 "100011111100000101111010",
						 "100011111100111100111111",
						 "100011111100111001010100",
						 "100011111100110101101001",
						 "100011111100110001111110",
						 "100011111100101110010011",
						 "100011111100101010101000",
						 "100011111100100110111101",
						 "100011111100100011010010",
						 "100011111100011111100111",
						 "100011111100011011111100",
						 "100011111100011000010001",
						 "100011111100010100100110",
						 "100011111100010000111011",
						 "100011111100001101010000",
						 "100011111100001001100101",
						 "100011111100000101111010",
						 "100011111100111100111111",
						 "100011111100111001010100",
						 "100011111100110101101001",
						 "100011111100110001111110",
						 "100011111100101110010011",
						 "100011111100101010101000",
						 "100011111100100110111101",
						 "100011111100100011010010",
						 "100011111100011111100111",
						 "100011111100011011111100",
						 "100011111100011000010001",
						 "100011111100010100100110",
						 "100011111100010000111011",
						 "100011111100001101010000",
						 "100011111100001001100101",
						 "100011111100000101111010",
						 "100011111010011010000001",
						 "100011111010010110010110",
						 "100011111010010010101011",
						 "100011111010001111000000",
						 "100011111010001011010101",
						 "100011111010000111101010",
						 "100011111010000011111111",
						 "100011111010000000010100",
						 "100011111001111100101001",
						 "100011111001111000111110",
						 "100011111001110101010011",
						 "100011111001110001101000",
						 "100011111001101101111101",
						 "100011111001101010010010",
						 "100011111001100110100111",
						 "100011111001100010111100",
						 "100011111010011010000001",
						 "100011111010010110010110",
						 "100011111010010010101011",
						 "100011111010001111000000",
						 "100011111010001011010101",
						 "100011111010000111101010",
						 "100011111010000011111111",
						 "100011111010000000010100",
						 "100011111001111100101001",
						 "100011111001111000111110",
						 "100011111001110101010011",
						 "100011111001110001101000",
						 "100011111001101101111101",
						 "100011111001101010010010",
						 "100011111001100110100111",
						 "100011111001100010111100",
						 "100011111010011010010000",
						 "100011111010010110100100",
						 "100011111010010010111000",
						 "100011111010001111001100",
						 "100011111010001011100000",
						 "100011111010000111110100",
						 "100011111010000100001000",
						 "100011111010000000011100",
						 "100011111001111100110000",
						 "100011111001111001000100",
						 "100011111001110101011000",
						 "100011111001110001101100",
						 "100011111001101110000000",
						 "100011111001101010010100",
						 "100011111001100110101000",
						 "100011111001100010111100",
						 "100011110111110111010010",
						 "100011110111110011100110",
						 "100011110111101111111010",
						 "100011110111101100001110",
						 "100011110111101000100010",
						 "100011110111100100110110",
						 "100011110111100001001010",
						 "100011110111011101011110",
						 "100011110111011001110010",
						 "100011110111010110000110",
						 "100011110111010010011010",
						 "100011110111001110101110",
						 "100011110111001011000010",
						 "100011110111000111010110",
						 "100011110111000011101010",
						 "100011110110111111111110",
						 "100011110111110111010010",
						 "100011110111110011100110",
						 "100011110111101111111010",
						 "100011110111101100001110",
						 "100011110111101000100010",
						 "100011110111100100110110",
						 "100011110111100001001010",
						 "100011110111011101011110",
						 "100011110111011001110010",
						 "100011110111010110000110",
						 "100011110111010010011010",
						 "100011110111001110101110",
						 "100011110111001011000010",
						 "100011110111000111010110",
						 "100011110111000011101010",
						 "100011110110111111111110",
						 "100011110111110111010010",
						 "100011110111110011100110",
						 "100011110111101111111010",
						 "100011110111101100001110",
						 "100011110111101000100010",
						 "100011110111100100110110",
						 "100011110111100001001010",
						 "100011110111011101011110",
						 "100011110111011001110010",
						 "100011110111010110000110",
						 "100011110111010010011010",
						 "100011110111001110101110",
						 "100011110111001011000010",
						 "100011110111000111010110",
						 "100011110111000011101010",
						 "100011110110111111111110",
						 "100011110101010100010100",
						 "100011110101010000101000",
						 "100011110101001100111100",
						 "100011110101001001010000",
						 "100011110101000101100100",
						 "100011110101000001111000",
						 "100011110100111110001100",
						 "100011110100111010100000",
						 "100011110100110110110100",
						 "100011110100110011001000",
						 "100011110100101111011100",
						 "100011110100101011110000",
						 "100011110100101000000100",
						 "100011110100100100011000",
						 "100011110100100000101100",
						 "100011110100011101000000",
						 "100011110101010100010100",
						 "100011110101010000101000",
						 "100011110101001100111100",
						 "100011110101001001010000",
						 "100011110101000101100100",
						 "100011110101000001111000",
						 "100011110100111110001100",
						 "100011110100111010100000",
						 "100011110100110110110100",
						 "100011110100110011001000",
						 "100011110100101111011100",
						 "100011110100101011110000",
						 "100011110100101000000100",
						 "100011110100100100011000",
						 "100011110100100000101100",
						 "100011110100011101000000",
						 "100011110010110001010110",
						 "100011110010101101101010",
						 "100011110010101001111110",
						 "100011110010100110010010",
						 "100011110010100010100110",
						 "100011110010011110111010",
						 "100011110010011011001110",
						 "100011110010010111100010",
						 "100011110010010011110110",
						 "100011110010010000001010",
						 "100011110010001100011110",
						 "100011110010001000110010",
						 "100011110010000101000110",
						 "100011110010000001011010",
						 "100011110001111101101110",
						 "100011110001111010000010",
						 "100011110010110001100101",
						 "100011110010101101111000",
						 "100011110010101010001011",
						 "100011110010100110011110",
						 "100011110010100010110001",
						 "100011110010011111000100",
						 "100011110010011011010111",
						 "100011110010010111101010",
						 "100011110010010011111101",
						 "100011110010010000010000",
						 "100011110010001100100011",
						 "100011110010001000110110",
						 "100011110010000101001001",
						 "100011110010000001011100",
						 "100011110001111101101111",
						 "100011110001111010000010",
						 "100011110010110001100101",
						 "100011110010101101111000",
						 "100011110010101010001011",
						 "100011110010100110011110",
						 "100011110010100010110001",
						 "100011110010011111000100",
						 "100011110010011011010111",
						 "100011110010010111101010",
						 "100011110010010011111101",
						 "100011110010010000010000",
						 "100011110010001100100011",
						 "100011110010001000110110",
						 "100011110010000101001001",
						 "100011110010000001011100",
						 "100011110001111101101111",
						 "100011110001111010000010",
						 "100011110000001110100111",
						 "100011110000001010111010",
						 "100011110000000111001101",
						 "100011110000000011100000",
						 "100011101111111111110011",
						 "100011101111111100000110",
						 "100011101111111000011001",
						 "100011101111110100101100",
						 "100011101111110000111111",
						 "100011101111101101010010",
						 "100011101111101001100101",
						 "100011101111100101111000",
						 "100011101111100010001011",
						 "100011101111011110011110",
						 "100011101111011010110001",
						 "100011101111010111000100",
						 "100011110000001110100111",
						 "100011110000001010111010",
						 "100011110000000111001101",
						 "100011110000000011100000",
						 "100011101111111111110011",
						 "100011101111111100000110",
						 "100011101111111000011001",
						 "100011101111110100101100",
						 "100011101111110000111111",
						 "100011101111101101010010",
						 "100011101111101001100101",
						 "100011101111100101111000",
						 "100011101111100010001011",
						 "100011101111011110011110",
						 "100011101111011010110001",
						 "100011101111010111000100",
						 "100011110000001110100111",
						 "100011110000001010111010",
						 "100011110000000111001101",
						 "100011110000000011100000",
						 "100011101111111111110011",
						 "100011101111111100000110",
						 "100011101111111000011001",
						 "100011101111110100101100",
						 "100011101111110000111111",
						 "100011101111101101010010",
						 "100011101111101001100101",
						 "100011101111100101111000",
						 "100011101111100010001011",
						 "100011101111011110011110",
						 "100011101111011010110001",
						 "100011101111010111000100",
						 "100011101101101011101001",
						 "100011101101100111111100",
						 "100011101101100100001111",
						 "100011101101100000100010",
						 "100011101101011100110101",
						 "100011101101011001001000",
						 "100011101101010101011011",
						 "100011101101010001101110",
						 "100011101101001110000001",
						 "100011101101001010010100",
						 "100011101101000110100111",
						 "100011101101000010111010",
						 "100011101100111111001101",
						 "100011101100111011100000",
						 "100011101100110111110011",
						 "100011101100110100000110",
						 "100011101101101011101001",
						 "100011101101100111111100",
						 "100011101101100100001111",
						 "100011101101100000100010",
						 "100011101101011100110101",
						 "100011101101011001001000",
						 "100011101101010101011011",
						 "100011101101010001101110",
						 "100011101101001110000001",
						 "100011101101001010010100",
						 "100011101101000110100111",
						 "100011101101000010111010",
						 "100011101100111111001101",
						 "100011101100111011100000",
						 "100011101100110111110011",
						 "100011101100110100000110",
						 "100011101101101011111000",
						 "100011101101101000001010",
						 "100011101101100100011100",
						 "100011101101100000101110",
						 "100011101101011101000000",
						 "100011101101011001010010",
						 "100011101101010101100100",
						 "100011101101010001110110",
						 "100011101101001110001000",
						 "100011101101001010011010",
						 "100011101101000110101100",
						 "100011101101000010111110",
						 "100011101100111111010000",
						 "100011101100111011100010",
						 "100011101100110111110100",
						 "100011101100110100000110",
						 "100011101011001000111010",
						 "100011101011000101001100",
						 "100011101011000001011110",
						 "100011101010111101110000",
						 "100011101010111010000010",
						 "100011101010110110010100",
						 "100011101010110010100110",
						 "100011101010101110111000",
						 "100011101010101011001010",
						 "100011101010100111011100",
						 "100011101010100011101110",
						 "100011101010100000000000",
						 "100011101010011100010010",
						 "100011101010011000100100",
						 "100011101010010100110110",
						 "100011101010010001001000",
						 "100011101011001000111010",
						 "100011101011000101001100",
						 "100011101011000001011110",
						 "100011101010111101110000",
						 "100011101010111010000010",
						 "100011101010110110010100",
						 "100011101010110010100110",
						 "100011101010101110111000",
						 "100011101010101011001010",
						 "100011101010100111011100",
						 "100011101010100011101110",
						 "100011101010100000000000",
						 "100011101010011100010010",
						 "100011101010011000100100",
						 "100011101010010100110110",
						 "100011101010010001001000",
						 "100011101000100101111100",
						 "100011101000100010001110",
						 "100011101000011110100000",
						 "100011101000011010110010",
						 "100011101000010111000100",
						 "100011101000010011010110",
						 "100011101000001111101000",
						 "100011101000001011111010",
						 "100011101000001000001100",
						 "100011101000000100011110",
						 "100011101000000000110000",
						 "100011100111111101000010",
						 "100011100111111001010100",
						 "100011100111110101100110",
						 "100011100111110001111000",
						 "100011100111101110001010",
						 "100011101000100101111100",
						 "100011101000100010001110",
						 "100011101000011110100000",
						 "100011101000011010110010",
						 "100011101000010111000100",
						 "100011101000010011010110",
						 "100011101000001111101000",
						 "100011101000001011111010",
						 "100011101000001000001100",
						 "100011101000000100011110",
						 "100011101000000000110000",
						 "100011100111111101000010",
						 "100011100111111001010100",
						 "100011100111110101100110",
						 "100011100111110001111000",
						 "100011100111101110001010",
						 "100011101000100101111100",
						 "100011101000100010001110",
						 "100011101000011110100000",
						 "100011101000011010110010",
						 "100011101000010111000100",
						 "100011101000010011010110",
						 "100011101000001111101000",
						 "100011101000001011111010",
						 "100011101000001000001100",
						 "100011101000000100011110",
						 "100011101000000000110000",
						 "100011100111111101000010",
						 "100011100111111001010100",
						 "100011100111110101100110",
						 "100011100111110001111000",
						 "100011100111101110001010",
						 "100011100110000010111110",
						 "100011100101111111010000",
						 "100011100101111011100010",
						 "100011100101110111110100",
						 "100011100101110100000110",
						 "100011100101110000011000",
						 "100011100101101100101010",
						 "100011100101101000111100",
						 "100011100101100101001110",
						 "100011100101100001100000",
						 "100011100101011101110010",
						 "100011100101011010000100",
						 "100011100101010110010110",
						 "100011100101010010101000",
						 "100011100101001110111010",
						 "100011100101001011001100",
						 "100011100110000011001101",
						 "100011100101111111011110",
						 "100011100101111011101111",
						 "100011100101111000000000",
						 "100011100101110100010001",
						 "100011100101110000100010",
						 "100011100101101100110011",
						 "100011100101101001000100",
						 "100011100101100101010101",
						 "100011100101100001100110",
						 "100011100101011101110111",
						 "100011100101011010001000",
						 "100011100101010110011001",
						 "100011100101010010101010",
						 "100011100101001110111011",
						 "100011100101001011001100",
						 "100011100110000011001101",
						 "100011100101111111011110",
						 "100011100101111011101111",
						 "100011100101111000000000",
						 "100011100101110100010001",
						 "100011100101110000100010",
						 "100011100101101100110011",
						 "100011100101101001000100",
						 "100011100101100101010101",
						 "100011100101100001100110",
						 "100011100101011101110111",
						 "100011100101011010001000",
						 "100011100101010110011001",
						 "100011100101010010101010",
						 "100011100101001110111011",
						 "100011100101001011001100",
						 "100011100011100000001111",
						 "100011100011011100100000",
						 "100011100011011000110001",
						 "100011100011010101000010",
						 "100011100011010001010011",
						 "100011100011001101100100",
						 "100011100011001001110101",
						 "100011100011000110000110",
						 "100011100011000010010111",
						 "100011100010111110101000",
						 "100011100010111010111001",
						 "100011100010110111001010",
						 "100011100010110011011011",
						 "100011100010101111101100",
						 "100011100010101011111101",
						 "100011100010101000001110",
						 "100011100011100000001111",
						 "100011100011011100100000",
						 "100011100011011000110001",
						 "100011100011010101000010",
						 "100011100011010001010011",
						 "100011100011001101100100",
						 "100011100011001001110101",
						 "100011100011000110000110",
						 "100011100011000010010111",
						 "100011100010111110101000",
						 "100011100010111010111001",
						 "100011100010110111001010",
						 "100011100010110011011011",
						 "100011100010101111101100",
						 "100011100010101011111101",
						 "100011100010101000001110",
						 "100011100000111101010001",
						 "100011100000111001100010",
						 "100011100000110101110011",
						 "100011100000110010000100",
						 "100011100000101110010101",
						 "100011100000101010100110",
						 "100011100000100110110111",
						 "100011100000100011001000",
						 "100011100000011111011001",
						 "100011100000011011101010",
						 "100011100000010111111011",
						 "100011100000010100001100",
						 "100011100000010000011101",
						 "100011100000001100101110",
						 "100011100000001000111111",
						 "100011100000000101010000",
						 "100011100000111101010001",
						 "100011100000111001100010",
						 "100011100000110101110011",
						 "100011100000110010000100",
						 "100011100000101110010101",
						 "100011100000101010100110",
						 "100011100000100110110111",
						 "100011100000100011001000",
						 "100011100000011111011001",
						 "100011100000011011101010",
						 "100011100000010111111011",
						 "100011100000010100001100",
						 "100011100000010000011101",
						 "100011100000001100101110",
						 "100011100000001000111111",
						 "100011100000000101010000",
						 "100011100000111101010001",
						 "100011100000111001100010",
						 "100011100000110101110011",
						 "100011100000110010000100",
						 "100011100000101110010101",
						 "100011100000101010100110",
						 "100011100000100110110111",
						 "100011100000100011001000",
						 "100011100000011111011001",
						 "100011100000011011101010",
						 "100011100000010111111011",
						 "100011100000010100001100",
						 "100011100000010000011101",
						 "100011100000001100101110",
						 "100011100000001000111111",
						 "100011100000000101010000",
						 "100011011110011010010011",
						 "100011011110010110100100",
						 "100011011110010010110101",
						 "100011011110001111000110",
						 "100011011110001011010111",
						 "100011011110000111101000",
						 "100011011110000011111001",
						 "100011011110000000001010",
						 "100011011101111100011011",
						 "100011011101111000101100",
						 "100011011101110100111101",
						 "100011011101110001001110",
						 "100011011101101101011111",
						 "100011011101101001110000",
						 "100011011101100110000001",
						 "100011011101100010010010",
						 "100011011110011010100010",
						 "100011011110010110110010",
						 "100011011110010011000010",
						 "100011011110001111010010",
						 "100011011110001011100010",
						 "100011011110000111110010",
						 "100011011110000100000010",
						 "100011011110000000010010",
						 "100011011101111100100010",
						 "100011011101111000110010",
						 "100011011101110101000010",
						 "100011011101110001010010",
						 "100011011101101101100010",
						 "100011011101101001110010",
						 "100011011101100110000010",
						 "100011011101100010010010",
						 "100011011110011010100010",
						 "100011011110010110110010",
						 "100011011110010011000010",
						 "100011011110001111010010",
						 "100011011110001011100010",
						 "100011011110000111110010",
						 "100011011110000100000010",
						 "100011011110000000010010",
						 "100011011101111100100010",
						 "100011011101111000110010",
						 "100011011101110101000010",
						 "100011011101110001010010",
						 "100011011101101101100010",
						 "100011011101101001110010",
						 "100011011101100110000010",
						 "100011011101100010010010",
						 "100011011011110111100100",
						 "100011011011110011110100",
						 "100011011011110000000100",
						 "100011011011101100010100",
						 "100011011011101000100100",
						 "100011011011100100110100",
						 "100011011011100001000100",
						 "100011011011011101010100",
						 "100011011011011001100100",
						 "100011011011010101110100",
						 "100011011011010010000100",
						 "100011011011001110010100",
						 "100011011011001010100100",
						 "100011011011000110110100",
						 "100011011011000011000100",
						 "100011011010111111010100",
						 "100011011011110111100100",
						 "100011011011110011110100",
						 "100011011011110000000100",
						 "100011011011101100010100",
						 "100011011011101000100100",
						 "100011011011100100110100",
						 "100011011011100001000100",
						 "100011011011011101010100",
						 "100011011011011001100100",
						 "100011011011010101110100",
						 "100011011011010010000100",
						 "100011011011001110010100",
						 "100011011011001010100100",
						 "100011011011000110110100",
						 "100011011011000011000100",
						 "100011011010111111010100",
						 "100011011011110111100100",
						 "100011011011110011110100",
						 "100011011011110000000100",
						 "100011011011101100010100",
						 "100011011011101000100100",
						 "100011011011100100110100",
						 "100011011011100001000100",
						 "100011011011011101010100",
						 "100011011011011001100100",
						 "100011011011010101110100",
						 "100011011011010010000100",
						 "100011011011001110010100",
						 "100011011011001010100100",
						 "100011011011000110110100",
						 "100011011011000011000100",
						 "100011011010111111010100",
						 "100011011001010100100110",
						 "100011011001010000110110",
						 "100011011001001101000110",
						 "100011011001001001010110",
						 "100011011001000101100110",
						 "100011011001000001110110",
						 "100011011000111110000110",
						 "100011011000111010010110",
						 "100011011000110110100110",
						 "100011011000110010110110",
						 "100011011000101111000110",
						 "100011011000101011010110",
						 "100011011000100111100110",
						 "100011011000100011110110",
						 "100011011000100000000110",
						 "100011011000011100010110",
						 "100011011001010100100110",
						 "100011011001010000110110",
						 "100011011001001101000110",
						 "100011011001001001010110",
						 "100011011001000101100110",
						 "100011011001000001110110",
						 "100011011000111110000110",
						 "100011011000111010010110",
						 "100011011000110110100110",
						 "100011011000110010110110",
						 "100011011000101111000110",
						 "100011011000101011010110",
						 "100011011000100111100110",
						 "100011011000100011110110",
						 "100011011000100000000110",
						 "100011011000011100010110",
						 "100011010110110001110111",
						 "100011010110101110000110",
						 "100011010110101010010101",
						 "100011010110100110100100",
						 "100011010110100010110011",
						 "100011010110011111000010",
						 "100011010110011011010001",
						 "100011010110010111100000",
						 "100011010110010011101111",
						 "100011010110001111111110",
						 "100011010110001100001101",
						 "100011010110001000011100",
						 "100011010110000100101011",
						 "100011010110000000111010",
						 "100011010101111101001001",
						 "100011010101111001011000",
						 "100011010110110001110111",
						 "100011010110101110000110",
						 "100011010110101010010101",
						 "100011010110100110100100",
						 "100011010110100010110011",
						 "100011010110011111000010",
						 "100011010110011011010001",
						 "100011010110010111100000",
						 "100011010110010011101111",
						 "100011010110001111111110",
						 "100011010110001100001101",
						 "100011010110001000011100",
						 "100011010110000100101011",
						 "100011010110000000111010",
						 "100011010101111101001001",
						 "100011010101111001011000",
						 "100011010110110001110111",
						 "100011010110101110000110",
						 "100011010110101010010101",
						 "100011010110100110100100",
						 "100011010110100010110011",
						 "100011010110011111000010",
						 "100011010110011011010001",
						 "100011010110010111100000",
						 "100011010110010011101111",
						 "100011010110001111111110",
						 "100011010110001100001101",
						 "100011010110001000011100",
						 "100011010110000100101011",
						 "100011010110000000111010",
						 "100011010101111101001001",
						 "100011010101111001011000",
						 "100011010100001110111001",
						 "100011010100001011001000",
						 "100011010100000111010111",
						 "100011010100000011100110",
						 "100011010011111111110101",
						 "100011010011111100000100",
						 "100011010011111000010011",
						 "100011010011110100100010",
						 "100011010011110000110001",
						 "100011010011101101000000",
						 "100011010011101001001111",
						 "100011010011100101011110",
						 "100011010011100001101101",
						 "100011010011011101111100",
						 "100011010011011010001011",
						 "100011010011010110011010",
						 "100011010100001110111001",
						 "100011010100001011001000",
						 "100011010100000111010111",
						 "100011010100000011100110",
						 "100011010011111111110101",
						 "100011010011111100000100",
						 "100011010011111000010011",
						 "100011010011110100100010",
						 "100011010011110000110001",
						 "100011010011101101000000",
						 "100011010011101001001111",
						 "100011010011100101011110",
						 "100011010011100001101101",
						 "100011010011011101111100",
						 "100011010011011010001011",
						 "100011010011010110011010",
						 "100011010100001110111001",
						 "100011010100001011001000",
						 "100011010100000111010111",
						 "100011010100000011100110",
						 "100011010011111111110101",
						 "100011010011111100000100",
						 "100011010011111000010011",
						 "100011010011110100100010",
						 "100011010011110000110001",
						 "100011010011101101000000",
						 "100011010011101001001111",
						 "100011010011100101011110",
						 "100011010011100001101101",
						 "100011010011011101111100",
						 "100011010011011010001011",
						 "100011010011010110011010",
						 "100011010001101011111011",
						 "100011010001101000001010",
						 "100011010001100100011001",
						 "100011010001100000101000",
						 "100011010001011100110111",
						 "100011010001011001000110",
						 "100011010001010101010101",
						 "100011010001010001100100",
						 "100011010001001101110011",
						 "100011010001001010000010",
						 "100011010001000110010001",
						 "100011010001000010100000",
						 "100011010000111110101111",
						 "100011010000111010111110",
						 "100011010000110111001101",
						 "100011010000110011011100",
						 "100011010001101011111011",
						 "100011010001101000001010",
						 "100011010001100100011001",
						 "100011010001100000101000",
						 "100011010001011100110111",
						 "100011010001011001000110",
						 "100011010001010101010101",
						 "100011010001010001100100",
						 "100011010001001101110011",
						 "100011010001001010000010",
						 "100011010001000110010001",
						 "100011010001000010100000",
						 "100011010000111110101111",
						 "100011010000111010111110",
						 "100011010000110111001101",
						 "100011010000110011011100",
						 "100011001111001001001100",
						 "100011001111000101011010",
						 "100011001111000001101000",
						 "100011001110111101110110",
						 "100011001110111010000100",
						 "100011001110110110010010",
						 "100011001110110010100000",
						 "100011001110101110101110",
						 "100011001110101010111100",
						 "100011001110100111001010",
						 "100011001110100011011000",
						 "100011001110011111100110",
						 "100011001110011011110100",
						 "100011001110011000000010",
						 "100011001110010100010000",
						 "100011001110010000011110",
						 "100011001111001001001100",
						 "100011001111000101011010",
						 "100011001111000001101000",
						 "100011001110111101110110",
						 "100011001110111010000100",
						 "100011001110110110010010",
						 "100011001110110010100000",
						 "100011001110101110101110",
						 "100011001110101010111100",
						 "100011001110100111001010",
						 "100011001110100011011000",
						 "100011001110011111100110",
						 "100011001110011011110100",
						 "100011001110011000000010",
						 "100011001110010100010000",
						 "100011001110010000011110",
						 "100011001111001001001100",
						 "100011001111000101011010",
						 "100011001111000001101000",
						 "100011001110111101110110",
						 "100011001110111010000100",
						 "100011001110110110010010",
						 "100011001110110010100000",
						 "100011001110101110101110",
						 "100011001110101010111100",
						 "100011001110100111001010",
						 "100011001110100011011000",
						 "100011001110011111100110",
						 "100011001110011011110100",
						 "100011001110011000000010",
						 "100011001110010100010000",
						 "100011001110010000011110",
						 "100011001100100110001110",
						 "100011001100100010011100",
						 "100011001100011110101010",
						 "100011001100011010111000",
						 "100011001100010111000110",
						 "100011001100010011010100",
						 "100011001100001111100010",
						 "100011001100001011110000",
						 "100011001100000111111110",
						 "100011001100000100001100",
						 "100011001100000000011010",
						 "100011001011111100101000",
						 "100011001011111000110110",
						 "100011001011110101000100",
						 "100011001011110001010010",
						 "100011001011101101100000",
						 "100011001100100110001110",
						 "100011001100100010011100",
						 "100011001100011110101010",
						 "100011001100011010111000",
						 "100011001100010111000110",
						 "100011001100010011010100",
						 "100011001100001111100010",
						 "100011001100001011110000",
						 "100011001100000111111110",
						 "100011001100000100001100",
						 "100011001100000000011010",
						 "100011001011111100101000",
						 "100011001011111000110110",
						 "100011001011110101000100",
						 "100011001011110001010010",
						 "100011001011101101100000",
						 "100011001100100110001110",
						 "100011001100100010011100",
						 "100011001100011110101010",
						 "100011001100011010111000",
						 "100011001100010111000110",
						 "100011001100010011010100",
						 "100011001100001111100010",
						 "100011001100001011110000",
						 "100011001100000111111110",
						 "100011001100000100001100",
						 "100011001100000000011010",
						 "100011001011111100101000",
						 "100011001011111000110110",
						 "100011001011110101000100",
						 "100011001011110001010010",
						 "100011001011101101100000",
						 "100011001010000011010000",
						 "100011001001111111011110",
						 "100011001001111011101100",
						 "100011001001110111111010",
						 "100011001001110100001000",
						 "100011001001110000010110",
						 "100011001001101100100100",
						 "100011001001101000110010",
						 "100011001001100101000000",
						 "100011001001100001001110",
						 "100011001001011101011100",
						 "100011001001011001101010",
						 "100011001001010101111000",
						 "100011001001010010000110",
						 "100011001001001110010100",
						 "100011001001001010100010",
						 "100011001010000011010000",
						 "100011001001111111011110",
						 "100011001001111011101100",
						 "100011001001110111111010",
						 "100011001001110100001000",
						 "100011001001110000010110",
						 "100011001001101100100100",
						 "100011001001101000110010",
						 "100011001001100101000000",
						 "100011001001100001001110",
						 "100011001001011101011100",
						 "100011001001011001101010",
						 "100011001001010101111000",
						 "100011001001010010000110",
						 "100011001001001110010100",
						 "100011001001001010100010",
						 "100011001010000011011111",
						 "100011001001111111101100",
						 "100011001001111011111001",
						 "100011001001111000000110",
						 "100011001001110100010011",
						 "100011001001110000100000",
						 "100011001001101100101101",
						 "100011001001101000111010",
						 "100011001001100101000111",
						 "100011001001100001010100",
						 "100011001001011101100001",
						 "100011001001011001101110",
						 "100011001001010101111011",
						 "100011001001010010001000",
						 "100011001001001110010101",
						 "100011001001001010100010",
						 "100011000111100000100001",
						 "100011000111011100101110",
						 "100011000111011000111011",
						 "100011000111010101001000",
						 "100011000111010001010101",
						 "100011000111001101100010",
						 "100011000111001001101111",
						 "100011000111000101111100",
						 "100011000111000010001001",
						 "100011000110111110010110",
						 "100011000110111010100011",
						 "100011000110110110110000",
						 "100011000110110010111101",
						 "100011000110101111001010",
						 "100011000110101011010111",
						 "100011000110100111100100",
						 "100011000111100000100001",
						 "100011000111011100101110",
						 "100011000111011000111011",
						 "100011000111010101001000",
						 "100011000111010001010101",
						 "100011000111001101100010",
						 "100011000111001001101111",
						 "100011000111000101111100",
						 "100011000111000010001001",
						 "100011000110111110010110",
						 "100011000110111010100011",
						 "100011000110110110110000",
						 "100011000110110010111101",
						 "100011000110101111001010",
						 "100011000110101011010111",
						 "100011000110100111100100",
						 "100011000100111101100011",
						 "100011000100111001110000",
						 "100011000100110101111101",
						 "100011000100110010001010",
						 "100011000100101110010111",
						 "100011000100101010100100",
						 "100011000100100110110001",
						 "100011000100100010111110",
						 "100011000100011111001011",
						 "100011000100011011011000",
						 "100011000100010111100101",
						 "100011000100010011110010",
						 "100011000100001111111111",
						 "100011000100001100001100",
						 "100011000100001000011001",
						 "100011000100000100100110",
						 "100011000100111101100011",
						 "100011000100111001110000",
						 "100011000100110101111101",
						 "100011000100110010001010",
						 "100011000100101110010111",
						 "100011000100101010100100",
						 "100011000100100110110001",
						 "100011000100100010111110",
						 "100011000100011111001011",
						 "100011000100011011011000",
						 "100011000100010111100101",
						 "100011000100010011110010",
						 "100011000100001111111111",
						 "100011000100001100001100",
						 "100011000100001000011001",
						 "100011000100000100100110",
						 "100011000100111101100011",
						 "100011000100111001110000",
						 "100011000100110101111101",
						 "100011000100110010001010",
						 "100011000100101110010111",
						 "100011000100101010100100",
						 "100011000100100110110001",
						 "100011000100100010111110",
						 "100011000100011111001011",
						 "100011000100011011011000",
						 "100011000100010111100101",
						 "100011000100010011110010",
						 "100011000100001111111111",
						 "100011000100001100001100",
						 "100011000100001000011001",
						 "100011000100000100100110",
						 "100011000010011010100101",
						 "100011000010010110110010",
						 "100011000010010010111111",
						 "100011000010001111001100",
						 "100011000010001011011001",
						 "100011000010000111100110",
						 "100011000010000011110011",
						 "100011000010000000000000",
						 "100011000001111100001101",
						 "100011000001111000011010",
						 "100011000001110100100111",
						 "100011000001110000110100",
						 "100011000001101101000001",
						 "100011000001101001001110",
						 "100011000001100101011011",
						 "100011000001100001101000",
						 "100011000010011010100101",
						 "100011000010010110110010",
						 "100011000010010010111111",
						 "100011000010001111001100",
						 "100011000010001011011001",
						 "100011000010000111100110",
						 "100011000010000011110011",
						 "100011000010000000000000",
						 "100011000001111100001101",
						 "100011000001111000011010",
						 "100011000001110100100111",
						 "100011000001110000110100",
						 "100011000001101101000001",
						 "100011000001101001001110",
						 "100011000001100101011011",
						 "100011000001100001101000",
						 "100011000010011010110100",
						 "100011000010010111000000",
						 "100011000010010011001100",
						 "100011000010001111011000",
						 "100011000010001011100100",
						 "100011000010000111110000",
						 "100011000010000011111100",
						 "100011000010000000001000",
						 "100011000001111100010100",
						 "100011000001111000100000",
						 "100011000001110100101100",
						 "100011000001110000111000",
						 "100011000001101101000100",
						 "100011000001101001010000",
						 "100011000001100101011100",
						 "100011000001100001101000",
						 "100010111111110111110110",
						 "100010111111110100000010",
						 "100010111111110000001110",
						 "100010111111101100011010",
						 "100010111111101000100110",
						 "100010111111100100110010",
						 "100010111111100000111110",
						 "100010111111011101001010",
						 "100010111111011001010110",
						 "100010111111010101100010",
						 "100010111111010001101110",
						 "100010111111001101111010",
						 "100010111111001010000110",
						 "100010111111000110010010",
						 "100010111111000010011110",
						 "100010111110111110101010",
						 "100010111111110111110110",
						 "100010111111110100000010",
						 "100010111111110000001110",
						 "100010111111101100011010",
						 "100010111111101000100110",
						 "100010111111100100110010",
						 "100010111111100000111110",
						 "100010111111011101001010",
						 "100010111111011001010110",
						 "100010111111010101100010",
						 "100010111111010001101110",
						 "100010111111001101111010",
						 "100010111111001010000110",
						 "100010111111000110010010",
						 "100010111111000010011110",
						 "100010111110111110101010",
						 "100010111101010100111000",
						 "100010111101010001000100",
						 "100010111101001101010000",
						 "100010111101001001011100",
						 "100010111101000101101000",
						 "100010111101000001110100",
						 "100010111100111110000000",
						 "100010111100111010001100",
						 "100010111100110110011000",
						 "100010111100110010100100",
						 "100010111100101110110000",
						 "100010111100101010111100",
						 "100010111100100111001000",
						 "100010111100100011010100",
						 "100010111100011111100000",
						 "100010111100011011101100",
						 "100010111101010100111000",
						 "100010111101010001000100",
						 "100010111101001101010000",
						 "100010111101001001011100",
						 "100010111101000101101000",
						 "100010111101000001110100",
						 "100010111100111110000000",
						 "100010111100111010001100",
						 "100010111100110110011000",
						 "100010111100110010100100",
						 "100010111100101110110000",
						 "100010111100101010111100",
						 "100010111100100111001000",
						 "100010111100100011010100",
						 "100010111100011111100000",
						 "100010111100011011101100",
						 "100010111101010100111000",
						 "100010111101010001000100",
						 "100010111101001101010000",
						 "100010111101001001011100",
						 "100010111101000101101000",
						 "100010111101000001110100",
						 "100010111100111110000000",
						 "100010111100111010001100",
						 "100010111100110110011000",
						 "100010111100110010100100",
						 "100010111100101110110000",
						 "100010111100101010111100",
						 "100010111100100111001000",
						 "100010111100100011010100",
						 "100010111100011111100000",
						 "100010111100011011101100",
						 "100010111010110001111010",
						 "100010111010101110000110",
						 "100010111010101010010010",
						 "100010111010100110011110",
						 "100010111010100010101010",
						 "100010111010011110110110",
						 "100010111010011011000010",
						 "100010111010010111001110",
						 "100010111010010011011010",
						 "100010111010001111100110",
						 "100010111010001011110010",
						 "100010111010000111111110",
						 "100010111010000100001010",
						 "100010111010000000010110",
						 "100010111001111100100010",
						 "100010111001111000101110",
						 "100010111010110001111010",
						 "100010111010101110000110",
						 "100010111010101010010010",
						 "100010111010100110011110",
						 "100010111010100010101010",
						 "100010111010011110110110",
						 "100010111010011011000010",
						 "100010111010010111001110",
						 "100010111010010011011010",
						 "100010111010001111100110",
						 "100010111010001011110010",
						 "100010111010000111111110",
						 "100010111010000100001010",
						 "100010111010000000010110",
						 "100010111001111100100010",
						 "100010111001111000101110",
						 "100010111010110001111010",
						 "100010111010101110000110",
						 "100010111010101010010010",
						 "100010111010100110011110",
						 "100010111010100010101010",
						 "100010111010011110110110",
						 "100010111010011011000010",
						 "100010111010010111001110",
						 "100010111010010011011010",
						 "100010111010001111100110",
						 "100010111010001011110010",
						 "100010111010000111111110",
						 "100010111010000100001010",
						 "100010111010000000010110",
						 "100010111001111100100010",
						 "100010111001111000101110",
						 "100010111000001111001011",
						 "100010111000001011010110",
						 "100010111000000111100001",
						 "100010111000000011101100",
						 "100010110111111111110111",
						 "100010110111111100000010",
						 "100010110111111000001101",
						 "100010110111110100011000",
						 "100010110111110000100011",
						 "100010110111101100101110",
						 "100010110111101000111001",
						 "100010110111100101000100",
						 "100010110111100001001111",
						 "100010110111011101011010",
						 "100010110111011001100101",
						 "100010110111010101110000",
						 "100010111000001111001011",
						 "100010111000001011010110",
						 "100010111000000111100001",
						 "100010111000000011101100",
						 "100010110111111111110111",
						 "100010110111111100000010",
						 "100010110111111000001101",
						 "100010110111110100011000",
						 "100010110111110000100011",
						 "100010110111101100101110",
						 "100010110111101000111001",
						 "100010110111100101000100",
						 "100010110111100001001111",
						 "100010110111011101011010",
						 "100010110111011001100101",
						 "100010110111010101110000",
						 "100010110101101100001101",
						 "100010110101101000011000",
						 "100010110101100100100011",
						 "100010110101100000101110",
						 "100010110101011100111001",
						 "100010110101011001000100",
						 "100010110101010101001111",
						 "100010110101010001011010",
						 "100010110101001101100101",
						 "100010110101001001110000",
						 "100010110101000101111011",
						 "100010110101000010000110",
						 "100010110100111110010001",
						 "100010110100111010011100",
						 "100010110100110110100111",
						 "100010110100110010110010",
						 "100010110101101100001101",
						 "100010110101101000011000",
						 "100010110101100100100011",
						 "100010110101100000101110",
						 "100010110101011100111001",
						 "100010110101011001000100",
						 "100010110101010101001111",
						 "100010110101010001011010",
						 "100010110101001101100101",
						 "100010110101001001110000",
						 "100010110101000101111011",
						 "100010110101000010000110",
						 "100010110100111110010001",
						 "100010110100111010011100",
						 "100010110100110110100111",
						 "100010110100110010110010",
						 "100010110101101100001101",
						 "100010110101101000011000",
						 "100010110101100100100011",
						 "100010110101100000101110",
						 "100010110101011100111001",
						 "100010110101011001000100",
						 "100010110101010101001111",
						 "100010110101010001011010",
						 "100010110101001101100101",
						 "100010110101001001110000",
						 "100010110101000101111011",
						 "100010110101000010000110",
						 "100010110100111110010001",
						 "100010110100111010011100",
						 "100010110100110110100111",
						 "100010110100110010110010",
						 "100010110011001001001111",
						 "100010110011000101011010",
						 "100010110011000001100101",
						 "100010110010111101110000",
						 "100010110010111001111011",
						 "100010110010110110000110",
						 "100010110010110010010001",
						 "100010110010101110011100",
						 "100010110010101010100111",
						 "100010110010100110110010",
						 "100010110010100010111101",
						 "100010110010011111001000",
						 "100010110010011011010011",
						 "100010110010010111011110",
						 "100010110010010011101001",
						 "100010110010001111110100",
						 "100010110011001001001111",
						 "100010110011000101011010",
						 "100010110011000001100101",
						 "100010110010111101110000",
						 "100010110010111001111011",
						 "100010110010110110000110",
						 "100010110010110010010001",
						 "100010110010101110011100",
						 "100010110010101010100111",
						 "100010110010100110110010",
						 "100010110010100010111101",
						 "100010110010011111001000",
						 "100010110010011011010011",
						 "100010110010010111011110",
						 "100010110010010011101001",
						 "100010110010001111110100",
						 "100010110011001001001111",
						 "100010110011000101011010",
						 "100010110011000001100101",
						 "100010110010111101110000",
						 "100010110010111001111011",
						 "100010110010110110000110",
						 "100010110010110010010001",
						 "100010110010101110011100",
						 "100010110010101010100111",
						 "100010110010100110110010",
						 "100010110010100010111101",
						 "100010110010011111001000",
						 "100010110010011011010011",
						 "100010110010010111011110",
						 "100010110010010011101001",
						 "100010110010001111110100",
						 "100010110000100110010001",
						 "100010110000100010011100",
						 "100010110000011110100111",
						 "100010110000011010110010",
						 "100010110000010110111101",
						 "100010110000010011001000",
						 "100010110000001111010011",
						 "100010110000001011011110",
						 "100010110000000111101001",
						 "100010110000000011110100",
						 "100010101111111111111111",
						 "100010101111111100001010",
						 "100010101111111000010101",
						 "100010101111110100100000",
						 "100010101111110000101011",
						 "100010101111101100110110",
						 "100010110000100110010001",
						 "100010110000100010011100",
						 "100010110000011110100111",
						 "100010110000011010110010",
						 "100010110000010110111101",
						 "100010110000010011001000",
						 "100010110000001111010011",
						 "100010110000001011011110",
						 "100010110000000111101001",
						 "100010110000000011110100",
						 "100010101111111111111111",
						 "100010101111111100001010",
						 "100010101111111000010101",
						 "100010101111110100100000",
						 "100010101111110000101011",
						 "100010101111101100110110",
						 "100010101110000011100010",
						 "100010101101111111101100",
						 "100010101101111011110110",
						 "100010101101111000000000",
						 "100010101101110100001010",
						 "100010101101110000010100",
						 "100010101101101100011110",
						 "100010101101101000101000",
						 "100010101101100100110010",
						 "100010101101100000111100",
						 "100010101101011101000110",
						 "100010101101011001010000",
						 "100010101101010101011010",
						 "100010101101010001100100",
						 "100010101101001101101110",
						 "100010101101001001111000",
						 "100010101110000011100010",
						 "100010101101111111101100",
						 "100010101101111011110110",
						 "100010101101111000000000",
						 "100010101101110100001010",
						 "100010101101110000010100",
						 "100010101101101100011110",
						 "100010101101101000101000",
						 "100010101101100100110010",
						 "100010101101100000111100",
						 "100010101101011101000110",
						 "100010101101011001010000",
						 "100010101101010101011010",
						 "100010101101010001100100",
						 "100010101101001101101110",
						 "100010101101001001111000",
						 "100010101110000011100010",
						 "100010101101111111101100",
						 "100010101101111011110110",
						 "100010101101111000000000",
						 "100010101101110100001010",
						 "100010101101110000010100",
						 "100010101101101100011110",
						 "100010101101101000101000",
						 "100010101101100100110010",
						 "100010101101100000111100",
						 "100010101101011101000110",
						 "100010101101011001010000",
						 "100010101101010101011010",
						 "100010101101010001100100",
						 "100010101101001101101110",
						 "100010101101001001111000",
						 "100010101011100000100100",
						 "100010101011011100101110",
						 "100010101011011000111000",
						 "100010101011010101000010",
						 "100010101011010001001100",
						 "100010101011001101010110",
						 "100010101011001001100000",
						 "100010101011000101101010",
						 "100010101011000001110100",
						 "100010101010111101111110",
						 "100010101010111010001000",
						 "100010101010110110010010",
						 "100010101010110010011100",
						 "100010101010101110100110",
						 "100010101010101010110000",
						 "100010101010100110111010",
						 "100010101011100000100100",
						 "100010101011011100101110",
						 "100010101011011000111000",
						 "100010101011010101000010",
						 "100010101011010001001100",
						 "100010101011001101010110",
						 "100010101011001001100000",
						 "100010101011000101101010",
						 "100010101011000001110100",
						 "100010101010111101111110",
						 "100010101010111010001000",
						 "100010101010110110010010",
						 "100010101010110010011100",
						 "100010101010101110100110",
						 "100010101010101010110000",
						 "100010101010100110111010",
						 "100010101011100000100100",
						 "100010101011011100101110",
						 "100010101011011000111000",
						 "100010101011010101000010",
						 "100010101011010001001100",
						 "100010101011001101010110",
						 "100010101011001001100000",
						 "100010101011000101101010",
						 "100010101011000001110100",
						 "100010101010111101111110",
						 "100010101010111010001000",
						 "100010101010110110010010",
						 "100010101010110010011100",
						 "100010101010101110100110",
						 "100010101010101010110000",
						 "100010101010100110111010",
						 "100010101000111101100110",
						 "100010101000111001110000",
						 "100010101000110101111010",
						 "100010101000110010000100",
						 "100010101000101110001110",
						 "100010101000101010011000",
						 "100010101000100110100010",
						 "100010101000100010101100",
						 "100010101000011110110110",
						 "100010101000011011000000",
						 "100010101000010111001010",
						 "100010101000010011010100",
						 "100010101000001111011110",
						 "100010101000001011101000",
						 "100010101000000111110010",
						 "100010101000000011111100",
						 "100010101000111101100110",
						 "100010101000111001110000",
						 "100010101000110101111010",
						 "100010101000110010000100",
						 "100010101000101110001110",
						 "100010101000101010011000",
						 "100010101000100110100010",
						 "100010101000100010101100",
						 "100010101000011110110110",
						 "100010101000011011000000",
						 "100010101000010111001010",
						 "100010101000010011010100",
						 "100010101000001111011110",
						 "100010101000001011101000",
						 "100010101000000111110010",
						 "100010101000000011111100",
						 "100010100110011010101000",
						 "100010100110010110110010",
						 "100010100110010010111100",
						 "100010100110001111000110",
						 "100010100110001011010000",
						 "100010100110000111011010",
						 "100010100110000011100100",
						 "100010100101111111101110",
						 "100010100101111011111000",
						 "100010100101111000000010",
						 "100010100101110100001100",
						 "100010100101110000010110",
						 "100010100101101100100000",
						 "100010100101101000101010",
						 "100010100101100100110100",
						 "100010100101100000111110",
						 "100010100110011010110111",
						 "100010100110010111000000",
						 "100010100110010011001001",
						 "100010100110001111010010",
						 "100010100110001011011011",
						 "100010100110000111100100",
						 "100010100110000011101101",
						 "100010100101111111110110",
						 "100010100101111011111111",
						 "100010100101111000001000",
						 "100010100101110100010001",
						 "100010100101110000011010",
						 "100010100101101100100011",
						 "100010100101101000101100",
						 "100010100101100100110101",
						 "100010100101100000111110",
						 "100010100110011010110111",
						 "100010100110010111000000",
						 "100010100110010011001001",
						 "100010100110001111010010",
						 "100010100110001011011011",
						 "100010100110000111100100",
						 "100010100110000011101101",
						 "100010100101111111110110",
						 "100010100101111011111111",
						 "100010100101111000001000",
						 "100010100101110100010001",
						 "100010100101110000011010",
						 "100010100101101100100011",
						 "100010100101101000101100",
						 "100010100101100100110101",
						 "100010100101100000111110",
						 "100010100011110111111001",
						 "100010100011110100000010",
						 "100010100011110000001011",
						 "100010100011101100010100",
						 "100010100011101000011101",
						 "100010100011100100100110",
						 "100010100011100000101111",
						 "100010100011011100111000",
						 "100010100011011001000001",
						 "100010100011010101001010",
						 "100010100011010001010011",
						 "100010100011001101011100",
						 "100010100011001001100101",
						 "100010100011000101101110",
						 "100010100011000001110111",
						 "100010100010111110000000",
						 "100010100011110111111001",
						 "100010100011110100000010",
						 "100010100011110000001011",
						 "100010100011101100010100",
						 "100010100011101000011101",
						 "100010100011100100100110",
						 "100010100011100000101111",
						 "100010100011011100111000",
						 "100010100011011001000001",
						 "100010100011010101001010",
						 "100010100011010001010011",
						 "100010100011001101011100",
						 "100010100011001001100101",
						 "100010100011000101101110",
						 "100010100011000001110111",
						 "100010100010111110000000",
						 "100010100001010100111011",
						 "100010100001010001000100",
						 "100010100001001101001101",
						 "100010100001001001010110",
						 "100010100001000101011111",
						 "100010100001000001101000",
						 "100010100000111101110001",
						 "100010100000111001111010",
						 "100010100000110110000011",
						 "100010100000110010001100",
						 "100010100000101110010101",
						 "100010100000101010011110",
						 "100010100000100110100111",
						 "100010100000100010110000",
						 "100010100000011110111001",
						 "100010100000011011000010",
						 "100010100001010100111011",
						 "100010100001010001000100",
						 "100010100001001101001101",
						 "100010100001001001010110",
						 "100010100001000101011111",
						 "100010100001000001101000",
						 "100010100000111101110001",
						 "100010100000111001111010",
						 "100010100000110110000011",
						 "100010100000110010001100",
						 "100010100000101110010101",
						 "100010100000101010011110",
						 "100010100000100110100111",
						 "100010100000100010110000",
						 "100010100000011110111001",
						 "100010100000011011000010",
						 "100010100001010100111011",
						 "100010100001010001000100",
						 "100010100001001101001101",
						 "100010100001001001010110",
						 "100010100001000101011111",
						 "100010100001000001101000",
						 "100010100000111101110001",
						 "100010100000111001111010",
						 "100010100000110110000011",
						 "100010100000110010001100",
						 "100010100000101110010101",
						 "100010100000101010011110",
						 "100010100000100110100111",
						 "100010100000100010110000",
						 "100010100000011110111001",
						 "100010100000011011000010",
						 "100010011110110001111101",
						 "100010011110101110000110",
						 "100010011110101010001111",
						 "100010011110100110011000",
						 "100010011110100010100001",
						 "100010011110011110101010",
						 "100010011110011010110011",
						 "100010011110010110111100",
						 "100010011110010011000101",
						 "100010011110001111001110",
						 "100010011110001011010111",
						 "100010011110000111100000",
						 "100010011110000011101001",
						 "100010011101111111110010",
						 "100010011101111011111011",
						 "100010011101111000000100",
						 "100010011110110001111101",
						 "100010011110101110000110",
						 "100010011110101010001111",
						 "100010011110100110011000",
						 "100010011110100010100001",
						 "100010011110011110101010",
						 "100010011110011010110011",
						 "100010011110010110111100",
						 "100010011110010011000101",
						 "100010011110001111001110",
						 "100010011110001011010111",
						 "100010011110000111100000",
						 "100010011110000011101001",
						 "100010011101111111110010",
						 "100010011101111011111011",
						 "100010011101111000000100",
						 "100010011110110001111101",
						 "100010011110101110000110",
						 "100010011110101010001111",
						 "100010011110100110011000",
						 "100010011110100010100001",
						 "100010011110011110101010",
						 "100010011110011010110011",
						 "100010011110010110111100",
						 "100010011110010011000101",
						 "100010011110001111001110",
						 "100010011110001011010111",
						 "100010011110000111100000",
						 "100010011110000011101001",
						 "100010011101111111110010",
						 "100010011101111011111011",
						 "100010011101111000000100",
						 "100010011100001110111111",
						 "100010011100001011001000",
						 "100010011100000111010001",
						 "100010011100000011011010",
						 "100010011011111111100011",
						 "100010011011111011101100",
						 "100010011011110111110101",
						 "100010011011110011111110",
						 "100010011011110000000111",
						 "100010011011101100010000",
						 "100010011011101000011001",
						 "100010011011100100100010",
						 "100010011011100000101011",
						 "100010011011011100110100",
						 "100010011011011000111101",
						 "100010011011010101000110",
						 "100010011100001111001110",
						 "100010011100001011010110",
						 "100010011100000111011110",
						 "100010011100000011100110",
						 "100010011011111111101110",
						 "100010011011111011110110",
						 "100010011011110111111110",
						 "100010011011110100000110",
						 "100010011011110000001110",
						 "100010011011101100010110",
						 "100010011011101000011110",
						 "100010011011100100100110",
						 "100010011011100000101110",
						 "100010011011011100110110",
						 "100010011011011000111110",
						 "100010011011010101000110",
						 "100010011001101100010000",
						 "100010011001101000011000",
						 "100010011001100100100000",
						 "100010011001100000101000",
						 "100010011001011100110000",
						 "100010011001011000111000",
						 "100010011001010101000000",
						 "100010011001010001001000",
						 "100010011001001101010000",
						 "100010011001001001011000",
						 "100010011001000101100000",
						 "100010011001000001101000",
						 "100010011000111101110000",
						 "100010011000111001111000",
						 "100010011000110110000000",
						 "100010011000110010001000",
						 "100010011001101100010000",
						 "100010011001101000011000",
						 "100010011001100100100000",
						 "100010011001100000101000",
						 "100010011001011100110000",
						 "100010011001011000111000",
						 "100010011001010101000000",
						 "100010011001010001001000",
						 "100010011001001101010000",
						 "100010011001001001011000",
						 "100010011001000101100000",
						 "100010011001000001101000",
						 "100010011000111101110000",
						 "100010011000111001111000",
						 "100010011000110110000000",
						 "100010011000110010001000",
						 "100010011001101100010000",
						 "100010011001101000011000",
						 "100010011001100100100000",
						 "100010011001100000101000",
						 "100010011001011100110000",
						 "100010011001011000111000",
						 "100010011001010101000000",
						 "100010011001010001001000",
						 "100010011001001101010000",
						 "100010011001001001011000",
						 "100010011001000101100000",
						 "100010011001000001101000",
						 "100010011000111101110000",
						 "100010011000111001111000",
						 "100010011000110110000000",
						 "100010011000110010001000",
						 "100010010111001001010010",
						 "100010010111000101011010",
						 "100010010111000001100010",
						 "100010010110111101101010",
						 "100010010110111001110010",
						 "100010010110110101111010",
						 "100010010110110010000010",
						 "100010010110101110001010",
						 "100010010110101010010010",
						 "100010010110100110011010",
						 "100010010110100010100010",
						 "100010010110011110101010",
						 "100010010110011010110010",
						 "100010010110010110111010",
						 "100010010110010011000010",
						 "100010010110001111001010",
						 "100010010111001001010010",
						 "100010010111000101011010",
						 "100010010111000001100010",
						 "100010010110111101101010",
						 "100010010110111001110010",
						 "100010010110110101111010",
						 "100010010110110010000010",
						 "100010010110101110001010",
						 "100010010110101010010010",
						 "100010010110100110011010",
						 "100010010110100010100010",
						 "100010010110011110101010",
						 "100010010110011010110010",
						 "100010010110010110111010",
						 "100010010110010011000010",
						 "100010010110001111001010",
						 "100010010111001001010010",
						 "100010010111000101011010",
						 "100010010111000001100010",
						 "100010010110111101101010",
						 "100010010110111001110010",
						 "100010010110110101111010",
						 "100010010110110010000010",
						 "100010010110101110001010",
						 "100010010110101010010010",
						 "100010010110100110011010",
						 "100010010110100010100010",
						 "100010010110011110101010",
						 "100010010110011010110010",
						 "100010010110010110111010",
						 "100010010110010011000010",
						 "100010010110001111001010",
						 "100010010100100110010100",
						 "100010010100100010011100",
						 "100010010100011110100100",
						 "100010010100011010101100",
						 "100010010100010110110100",
						 "100010010100010010111100",
						 "100010010100001111000100",
						 "100010010100001011001100",
						 "100010010100000111010100",
						 "100010010100000011011100",
						 "100010010011111111100100",
						 "100010010011111011101100",
						 "100010010011110111110100",
						 "100010010011110011111100",
						 "100010010011110000000100",
						 "100010010011101100001100",
						 "100010010100100110010100",
						 "100010010100100010011100",
						 "100010010100011110100100",
						 "100010010100011010101100",
						 "100010010100010110110100",
						 "100010010100010010111100",
						 "100010010100001111000100",
						 "100010010100001011001100",
						 "100010010100000111010100",
						 "100010010100000011011100",
						 "100010010011111111100100",
						 "100010010011111011101100",
						 "100010010011110111110100",
						 "100010010011110011111100",
						 "100010010011110000000100",
						 "100010010011101100001100",
						 "100010010010000011010110",
						 "100010010001111111011110",
						 "100010010001111011100110",
						 "100010010001110111101110",
						 "100010010001110011110110",
						 "100010010001101111111110",
						 "100010010001101100000110",
						 "100010010001101000001110",
						 "100010010001100100010110",
						 "100010010001100000011110",
						 "100010010001011100100110",
						 "100010010001011000101110",
						 "100010010001010100110110",
						 "100010010001010000111110",
						 "100010010001001101000110",
						 "100010010001001001001110",
						 "100010010010000011100101",
						 "100010010001111111101100",
						 "100010010001111011110011",
						 "100010010001110111111010",
						 "100010010001110100000001",
						 "100010010001110000001000",
						 "100010010001101100001111",
						 "100010010001101000010110",
						 "100010010001100100011101",
						 "100010010001100000100100",
						 "100010010001011100101011",
						 "100010010001011000110010",
						 "100010010001010100111001",
						 "100010010001010001000000",
						 "100010010001001101000111",
						 "100010010001001001001110",
						 "100010010010000011100101",
						 "100010010001111111101100",
						 "100010010001111011110011",
						 "100010010001110111111010",
						 "100010010001110100000001",
						 "100010010001110000001000",
						 "100010010001101100001111",
						 "100010010001101000010110",
						 "100010010001100100011101",
						 "100010010001100000100100",
						 "100010010001011100101011",
						 "100010010001011000110010",
						 "100010010001010100111001",
						 "100010010001010001000000",
						 "100010010001001101000111",
						 "100010010001001001001110",
						 "100010001111100000100111",
						 "100010001111011100101110",
						 "100010001111011000110101",
						 "100010001111010100111100",
						 "100010001111010001000011",
						 "100010001111001101001010",
						 "100010001111001001010001",
						 "100010001111000101011000",
						 "100010001111000001011111",
						 "100010001110111101100110",
						 "100010001110111001101101",
						 "100010001110110101110100",
						 "100010001110110001111011",
						 "100010001110101110000010",
						 "100010001110101010001001",
						 "100010001110100110010000",
						 "100010001111100000100111",
						 "100010001111011100101110",
						 "100010001111011000110101",
						 "100010001111010100111100",
						 "100010001111010001000011",
						 "100010001111001101001010",
						 "100010001111001001010001",
						 "100010001111000101011000",
						 "100010001111000001011111",
						 "100010001110111101100110",
						 "100010001110111001101101",
						 "100010001110110101110100",
						 "100010001110110001111011",
						 "100010001110101110000010",
						 "100010001110101010001001",
						 "100010001110100110010000",
						 "100010001100111101101001",
						 "100010001100111001110000",
						 "100010001100110101110111",
						 "100010001100110001111110",
						 "100010001100101110000101",
						 "100010001100101010001100",
						 "100010001100100110010011",
						 "100010001100100010011010",
						 "100010001100011110100001",
						 "100010001100011010101000",
						 "100010001100010110101111",
						 "100010001100010010110110",
						 "100010001100001110111101",
						 "100010001100001011000100",
						 "100010001100000111001011",
						 "100010001100000011010010",
						 "100010001100111101101001",
						 "100010001100111001110000",
						 "100010001100110101110111",
						 "100010001100110001111110",
						 "100010001100101110000101",
						 "100010001100101010001100",
						 "100010001100100110010011",
						 "100010001100100010011010",
						 "100010001100011110100001",
						 "100010001100011010101000",
						 "100010001100010110101111",
						 "100010001100010010110110",
						 "100010001100001110111101",
						 "100010001100001011000100",
						 "100010001100000111001011",
						 "100010001100000011010010",
						 "100010001100111101101001",
						 "100010001100111001110000",
						 "100010001100110101110111",
						 "100010001100110001111110",
						 "100010001100101110000101",
						 "100010001100101010001100",
						 "100010001100100110010011",
						 "100010001100100010011010",
						 "100010001100011110100001",
						 "100010001100011010101000",
						 "100010001100010110101111",
						 "100010001100010010110110",
						 "100010001100001110111101",
						 "100010001100001011000100",
						 "100010001100000111001011",
						 "100010001100000011010010",
						 "100010001010011010101011",
						 "100010001010010110110010",
						 "100010001010010010111001",
						 "100010001010001111000000",
						 "100010001010001011000111",
						 "100010001010000111001110",
						 "100010001010000011010101",
						 "100010001001111111011100",
						 "100010001001111011100011",
						 "100010001001110111101010",
						 "100010001001110011110001",
						 "100010001001101111111000",
						 "100010001001101011111111",
						 "100010001001101000000110",
						 "100010001001100100001101",
						 "100010001001100000010100",
						 "100010001010011010101011",
						 "100010001010010110110010",
						 "100010001010010010111001",
						 "100010001010001111000000",
						 "100010001010001011000111",
						 "100010001010000111001110",
						 "100010001010000011010101",
						 "100010001001111111011100",
						 "100010001001111011100011",
						 "100010001001110111101010",
						 "100010001001110011110001",
						 "100010001001101111111000",
						 "100010001001101011111111",
						 "100010001001101000000110",
						 "100010001001100100001101",
						 "100010001001100000010100",
						 "100010001010011010101011",
						 "100010001010010110110010",
						 "100010001010010010111001",
						 "100010001010001111000000",
						 "100010001010001011000111",
						 "100010001010000111001110",
						 "100010001010000011010101",
						 "100010001001111111011100",
						 "100010001001111011100011",
						 "100010001001110111101010",
						 "100010001001110011110001",
						 "100010001001101111111000",
						 "100010001001101011111111",
						 "100010001001101000000110",
						 "100010001001100100001101",
						 "100010001001100000010100",
						 "100010000111110111101101",
						 "100010000111110011110100",
						 "100010000111101111111011",
						 "100010000111101100000010",
						 "100010000111101000001001",
						 "100010000111100100010000",
						 "100010000111100000010111",
						 "100010000111011100011110",
						 "100010000111011000100101",
						 "100010000111010100101100",
						 "100010000111010000110011",
						 "100010000111001100111010",
						 "100010000111001001000001",
						 "100010000111000101001000",
						 "100010000111000001001111",
						 "100010000110111101010110",
						 "100010000111110111101101",
						 "100010000111110011110100",
						 "100010000111101111111011",
						 "100010000111101100000010",
						 "100010000111101000001001",
						 "100010000111100100010000",
						 "100010000111100000010111",
						 "100010000111011100011110",
						 "100010000111011000100101",
						 "100010000111010100101100",
						 "100010000111010000110011",
						 "100010000111001100111010",
						 "100010000111001001000001",
						 "100010000111000101001000",
						 "100010000111000001001111",
						 "100010000110111101010110",
						 "100010000101010100111110",
						 "100010000101010001000100",
						 "100010000101001101001010",
						 "100010000101001001010000",
						 "100010000101000101010110",
						 "100010000101000001011100",
						 "100010000100111101100010",
						 "100010000100111001101000",
						 "100010000100110101101110",
						 "100010000100110001110100",
						 "100010000100101101111010",
						 "100010000100101010000000",
						 "100010000100100110000110",
						 "100010000100100010001100",
						 "100010000100011110010010",
						 "100010000100011010011000",
						 "100010000101010100111110",
						 "100010000101010001000100",
						 "100010000101001101001010",
						 "100010000101001001010000",
						 "100010000101000101010110",
						 "100010000101000001011100",
						 "100010000100111101100010",
						 "100010000100111001101000",
						 "100010000100110101101110",
						 "100010000100110001110100",
						 "100010000100101101111010",
						 "100010000100101010000000",
						 "100010000100100110000110",
						 "100010000100100010001100",
						 "100010000100011110010010",
						 "100010000100011010011000",
						 "100010000101010100111110",
						 "100010000101010001000100",
						 "100010000101001101001010",
						 "100010000101001001010000",
						 "100010000101000101010110",
						 "100010000101000001011100",
						 "100010000100111101100010",
						 "100010000100111001101000",
						 "100010000100110101101110",
						 "100010000100110001110100",
						 "100010000100101101111010",
						 "100010000100101010000000",
						 "100010000100100110000110",
						 "100010000100100010001100",
						 "100010000100011110010010",
						 "100010000100011010011000",
						 "100010000010110010000000",
						 "100010000010101110000110",
						 "100010000010101010001100",
						 "100010000010100110010010",
						 "100010000010100010011000",
						 "100010000010011110011110",
						 "100010000010011010100100",
						 "100010000010010110101010",
						 "100010000010010010110000",
						 "100010000010001110110110",
						 "100010000010001010111100",
						 "100010000010000111000010",
						 "100010000010000011001000",
						 "100010000001111111001110",
						 "100010000001111011010100",
						 "100010000001110111011010",
						 "100010000010110010000000",
						 "100010000010101110000110",
						 "100010000010101010001100",
						 "100010000010100110010010",
						 "100010000010100010011000",
						 "100010000010011110011110",
						 "100010000010011010100100",
						 "100010000010010110101010",
						 "100010000010010010110000",
						 "100010000010001110110110",
						 "100010000010001010111100",
						 "100010000010000111000010",
						 "100010000010000011001000",
						 "100010000001111111001110",
						 "100010000001111011010100",
						 "100010000001110111011010",
						 "100010000010110010000000",
						 "100010000010101110000110",
						 "100010000010101010001100",
						 "100010000010100110010010",
						 "100010000010100010011000",
						 "100010000010011110011110",
						 "100010000010011010100100",
						 "100010000010010110101010",
						 "100010000010010010110000",
						 "100010000010001110110110",
						 "100010000010001010111100",
						 "100010000010000111000010",
						 "100010000010000011001000",
						 "100010000001111111001110",
						 "100010000001111011010100",
						 "100010000001110111011010",
						 "100010000000001111000010",
						 "100010000000001011001000",
						 "100010000000000111001110",
						 "100010000000000011010100",
						 "100001111111111111011010",
						 "100001111111111011100000",
						 "100001111111110111100110",
						 "100001111111110011101100",
						 "100001111111101111110010",
						 "100001111111101011111000",
						 "100001111111100111111110",
						 "100001111111100100000100",
						 "100001111111100000001010",
						 "100001111111011100010000",
						 "100001111111011000010110",
						 "100001111111010100011100",
						 "100010000000001111000010",
						 "100010000000001011001000",
						 "100010000000000111001110",
						 "100010000000000011010100",
						 "100001111111111111011010",
						 "100001111111111011100000",
						 "100001111111110111100110",
						 "100001111111110011101100",
						 "100001111111101111110010",
						 "100001111111101011111000",
						 "100001111111100111111110",
						 "100001111111100100000100",
						 "100001111111100000001010",
						 "100001111111011100010000",
						 "100001111111011000010110",
						 "100001111111010100011100",
						 "100001111101101100000100",
						 "100001111101101000001010",
						 "100001111101100100010000",
						 "100001111101100000010110",
						 "100001111101011100011100",
						 "100001111101011000100010",
						 "100001111101010100101000",
						 "100001111101010000101110",
						 "100001111101001100110100",
						 "100001111101001000111010",
						 "100001111101000101000000",
						 "100001111101000001000110",
						 "100001111100111101001100",
						 "100001111100111001010010",
						 "100001111100110101011000",
						 "100001111100110001011110",
						 "100001111101101100000100",
						 "100001111101101000001010",
						 "100001111101100100010000",
						 "100001111101100000010110",
						 "100001111101011100011100",
						 "100001111101011000100010",
						 "100001111101010100101000",
						 "100001111101010000101110",
						 "100001111101001100110100",
						 "100001111101001000111010",
						 "100001111101000101000000",
						 "100001111101000001000110",
						 "100001111100111101001100",
						 "100001111100111001010010",
						 "100001111100110101011000",
						 "100001111100110001011110",
						 "100001111101101100000100",
						 "100001111101101000001010",
						 "100001111101100100010000",
						 "100001111101100000010110",
						 "100001111101011100011100",
						 "100001111101011000100010",
						 "100001111101010100101000",
						 "100001111101010000101110",
						 "100001111101001100110100",
						 "100001111101001000111010",
						 "100001111101000101000000",
						 "100001111101000001000110",
						 "100001111100111101001100",
						 "100001111100111001010010",
						 "100001111100110101011000",
						 "100001111100110001011110",
						 "100001111011001001000110",
						 "100001111011000101001100",
						 "100001111011000001010010",
						 "100001111010111101011000",
						 "100001111010111001011110",
						 "100001111010110101100100",
						 "100001111010110001101010",
						 "100001111010101101110000",
						 "100001111010101001110110",
						 "100001111010100101111100",
						 "100001111010100010000010",
						 "100001111010011110001000",
						 "100001111010011010001110",
						 "100001111010010110010100",
						 "100001111010010010011010",
						 "100001111010001110100000",
						 "100001111011001001000110",
						 "100001111011000101001100",
						 "100001111011000001010010",
						 "100001111010111101011000",
						 "100001111010111001011110",
						 "100001111010110101100100",
						 "100001111010110001101010",
						 "100001111010101101110000",
						 "100001111010101001110110",
						 "100001111010100101111100",
						 "100001111010100010000010",
						 "100001111010011110001000",
						 "100001111010011010001110",
						 "100001111010010110010100",
						 "100001111010010010011010",
						 "100001111010001110100000",
						 "100001111000100110010111",
						 "100001111000100010011100",
						 "100001111000011110100001",
						 "100001111000011010100110",
						 "100001111000010110101011",
						 "100001111000010010110000",
						 "100001111000001110110101",
						 "100001111000001010111010",
						 "100001111000000110111111",
						 "100001111000000011000100",
						 "100001110111111111001001",
						 "100001110111111011001110",
						 "100001110111110111010011",
						 "100001110111110011011000",
						 "100001110111101111011101",
						 "100001110111101011100010",
						 "100001111000100110010111",
						 "100001111000100010011100",
						 "100001111000011110100001",
						 "100001111000011010100110",
						 "100001111000010110101011",
						 "100001111000010010110000",
						 "100001111000001110110101",
						 "100001111000001010111010",
						 "100001111000000110111111",
						 "100001111000000011000100",
						 "100001110111111111001001",
						 "100001110111111011001110",
						 "100001110111110111010011",
						 "100001110111110011011000",
						 "100001110111101111011101",
						 "100001110111101011100010",
						 "100001111000100110010111",
						 "100001111000100010011100",
						 "100001111000011110100001",
						 "100001111000011010100110",
						 "100001111000010110101011",
						 "100001111000010010110000",
						 "100001111000001110110101",
						 "100001111000001010111010",
						 "100001111000000110111111",
						 "100001111000000011000100",
						 "100001110111111111001001",
						 "100001110111111011001110",
						 "100001110111110111010011",
						 "100001110111110011011000",
						 "100001110111101111011101",
						 "100001110111101011100010",
						 "100001110110000011011001",
						 "100001110101111111011110",
						 "100001110101111011100011",
						 "100001110101110111101000",
						 "100001110101110011101101",
						 "100001110101101111110010",
						 "100001110101101011110111",
						 "100001110101100111111100",
						 "100001110101100100000001",
						 "100001110101100000000110",
						 "100001110101011100001011",
						 "100001110101011000010000",
						 "100001110101010100010101",
						 "100001110101010000011010",
						 "100001110101001100011111",
						 "100001110101001000100100",
						 "100001110110000011011001",
						 "100001110101111111011110",
						 "100001110101111011100011",
						 "100001110101110111101000",
						 "100001110101110011101101",
						 "100001110101101111110010",
						 "100001110101101011110111",
						 "100001110101100111111100",
						 "100001110101100100000001",
						 "100001110101100000000110",
						 "100001110101011100001011",
						 "100001110101011000010000",
						 "100001110101010100010101",
						 "100001110101010000011010",
						 "100001110101001100011111",
						 "100001110101001000100100",
						 "100001110110000011011001",
						 "100001110101111111011110",
						 "100001110101111011100011",
						 "100001110101110111101000",
						 "100001110101110011101101",
						 "100001110101101111110010",
						 "100001110101101011110111",
						 "100001110101100111111100",
						 "100001110101100100000001",
						 "100001110101100000000110",
						 "100001110101011100001011",
						 "100001110101011000010000",
						 "100001110101010100010101",
						 "100001110101010000011010",
						 "100001110101001100011111",
						 "100001110101001000100100",
						 "100001110011100000011011",
						 "100001110011011100100000",
						 "100001110011011000100101",
						 "100001110011010100101010",
						 "100001110011010000101111",
						 "100001110011001100110100",
						 "100001110011001000111001",
						 "100001110011000100111110",
						 "100001110011000001000011",
						 "100001110010111101001000",
						 "100001110010111001001101",
						 "100001110010110101010010",
						 "100001110010110001010111",
						 "100001110010101101011100",
						 "100001110010101001100001",
						 "100001110010100101100110",
						 "100001110011100000011011",
						 "100001110011011100100000",
						 "100001110011011000100101",
						 "100001110011010100101010",
						 "100001110011010000101111",
						 "100001110011001100110100",
						 "100001110011001000111001",
						 "100001110011000100111110",
						 "100001110011000001000011",
						 "100001110010111101001000",
						 "100001110010111001001101",
						 "100001110010110101010010",
						 "100001110010110001010111",
						 "100001110010101101011100",
						 "100001110010101001100001",
						 "100001110010100101100110",
						 "100001110000111101011101",
						 "100001110000111001100010",
						 "100001110000110101100111",
						 "100001110000110001101100",
						 "100001110000101101110001",
						 "100001110000101001110110",
						 "100001110000100101111011",
						 "100001110000100010000000",
						 "100001110000011110000101",
						 "100001110000011010001010",
						 "100001110000010110001111",
						 "100001110000010010010100",
						 "100001110000001110011001",
						 "100001110000001010011110",
						 "100001110000000110100011",
						 "100001110000000010101000",
						 "100001110000111101011101",
						 "100001110000111001100010",
						 "100001110000110101100111",
						 "100001110000110001101100",
						 "100001110000101101110001",
						 "100001110000101001110110",
						 "100001110000100101111011",
						 "100001110000100010000000",
						 "100001110000011110000101",
						 "100001110000011010001010",
						 "100001110000010110001111",
						 "100001110000010010010100",
						 "100001110000001110011001",
						 "100001110000001010011110",
						 "100001110000000110100011",
						 "100001110000000010101000",
						 "100001110000111101011101",
						 "100001110000111001100010",
						 "100001110000110101100111",
						 "100001110000110001101100",
						 "100001110000101101110001",
						 "100001110000101001110110",
						 "100001110000100101111011",
						 "100001110000100010000000",
						 "100001110000011110000101",
						 "100001110000011010001010",
						 "100001110000010110001111",
						 "100001110000010010010100",
						 "100001110000001110011001",
						 "100001110000001010011110",
						 "100001110000000110100011",
						 "100001110000000010101000",
						 "100001101110011010011111",
						 "100001101110010110100100",
						 "100001101110010010101001",
						 "100001101110001110101110",
						 "100001101110001010110011",
						 "100001101110000110111000",
						 "100001101110000010111101",
						 "100001101101111111000010",
						 "100001101101111011000111",
						 "100001101101110111001100",
						 "100001101101110011010001",
						 "100001101101101111010110",
						 "100001101101101011011011",
						 "100001101101100111100000",
						 "100001101101100011100101",
						 "100001101101011111101010",
						 "100001101110011010011111",
						 "100001101110010110100100",
						 "100001101110010010101001",
						 "100001101110001110101110",
						 "100001101110001010110011",
						 "100001101110000110111000",
						 "100001101110000010111101",
						 "100001101101111111000010",
						 "100001101101111011000111",
						 "100001101101110111001100",
						 "100001101101110011010001",
						 "100001101101101111010110",
						 "100001101101101011011011",
						 "100001101101100111100000",
						 "100001101101100011100101",
						 "100001101101011111101010",
						 "100001101011110111100001",
						 "100001101011110011100110",
						 "100001101011101111101011",
						 "100001101011101011110000",
						 "100001101011100111110101",
						 "100001101011100011111010",
						 "100001101011011111111111",
						 "100001101011011100000100",
						 "100001101011011000001001",
						 "100001101011010100001110",
						 "100001101011010000010011",
						 "100001101011001100011000",
						 "100001101011001000011101",
						 "100001101011000100100010",
						 "100001101011000000100111",
						 "100001101010111100101100",
						 "100001101011110111100001",
						 "100001101011110011100110",
						 "100001101011101111101011",
						 "100001101011101011110000",
						 "100001101011100111110101",
						 "100001101011100011111010",
						 "100001101011011111111111",
						 "100001101011011100000100",
						 "100001101011011000001001",
						 "100001101011010100001110",
						 "100001101011010000010011",
						 "100001101011001100011000",
						 "100001101011001000011101",
						 "100001101011000100100010",
						 "100001101011000000100111",
						 "100001101010111100101100",
						 "100001101011110111110000",
						 "100001101011110011110100",
						 "100001101011101111111000",
						 "100001101011101011111100",
						 "100001101011101000000000",
						 "100001101011100100000100",
						 "100001101011100000001000",
						 "100001101011011100001100",
						 "100001101011011000010000",
						 "100001101011010100010100",
						 "100001101011010000011000",
						 "100001101011001100011100",
						 "100001101011001000100000",
						 "100001101011000100100100",
						 "100001101011000000101000",
						 "100001101010111100101100",
						 "100001101001010100110010",
						 "100001101001010000110110",
						 "100001101001001100111010",
						 "100001101001001000111110",
						 "100001101001000101000010",
						 "100001101001000001000110",
						 "100001101000111101001010",
						 "100001101000111001001110",
						 "100001101000110101010010",
						 "100001101000110001010110",
						 "100001101000101101011010",
						 "100001101000101001011110",
						 "100001101000100101100010",
						 "100001101000100001100110",
						 "100001101000011101101010",
						 "100001101000011001101110",
						 "100001101001010100110010",
						 "100001101001010000110110",
						 "100001101001001100111010",
						 "100001101001001000111110",
						 "100001101001000101000010",
						 "100001101001000001000110",
						 "100001101000111101001010",
						 "100001101000111001001110",
						 "100001101000110101010010",
						 "100001101000110001010110",
						 "100001101000101101011010",
						 "100001101000101001011110",
						 "100001101000100101100010",
						 "100001101000100001100110",
						 "100001101000011101101010",
						 "100001101000011001101110",
						 "100001101001010100110010",
						 "100001101001010000110110",
						 "100001101001001100111010",
						 "100001101001001000111110",
						 "100001101001000101000010",
						 "100001101001000001000110",
						 "100001101000111101001010",
						 "100001101000111001001110",
						 "100001101000110101010010",
						 "100001101000110001010110",
						 "100001101000101101011010",
						 "100001101000101001011110",
						 "100001101000100101100010",
						 "100001101000100001100110",
						 "100001101000011101101010",
						 "100001101000011001101110",
						 "100001100110110001110100",
						 "100001100110101101111000",
						 "100001100110101001111100",
						 "100001100110100110000000",
						 "100001100110100010000100",
						 "100001100110011110001000",
						 "100001100110011010001100",
						 "100001100110010110010000",
						 "100001100110010010010100",
						 "100001100110001110011000",
						 "100001100110001010011100",
						 "100001100110000110100000",
						 "100001100110000010100100",
						 "100001100101111110101000",
						 "100001100101111010101100",
						 "100001100101110110110000",
						 "100001100110110001110100",
						 "100001100110101101111000",
						 "100001100110101001111100",
						 "100001100110100110000000",
						 "100001100110100010000100",
						 "100001100110011110001000",
						 "100001100110011010001100",
						 "100001100110010110010000",
						 "100001100110010010010100",
						 "100001100110001110011000",
						 "100001100110001010011100",
						 "100001100110000110100000",
						 "100001100110000010100100",
						 "100001100101111110101000",
						 "100001100101111010101100",
						 "100001100101110110110000",
						 "100001100100001110110110",
						 "100001100100001010111010",
						 "100001100100000110111110",
						 "100001100100000011000010",
						 "100001100011111111000110",
						 "100001100011111011001010",
						 "100001100011110111001110",
						 "100001100011110011010010",
						 "100001100011101111010110",
						 "100001100011101011011010",
						 "100001100011100111011110",
						 "100001100011100011100010",
						 "100001100011011111100110",
						 "100001100011011011101010",
						 "100001100011010111101110",
						 "100001100011010011110010",
						 "100001100100001110110110",
						 "100001100100001010111010",
						 "100001100100000110111110",
						 "100001100100000011000010",
						 "100001100011111111000110",
						 "100001100011111011001010",
						 "100001100011110111001110",
						 "100001100011110011010010",
						 "100001100011101111010110",
						 "100001100011101011011010",
						 "100001100011100111011110",
						 "100001100011100011100010",
						 "100001100011011111100110",
						 "100001100011011011101010",
						 "100001100011010111101110",
						 "100001100011010011110010",
						 "100001100100001110110110",
						 "100001100100001010111010",
						 "100001100100000110111110",
						 "100001100100000011000010",
						 "100001100011111111000110",
						 "100001100011111011001010",
						 "100001100011110111001110",
						 "100001100011110011010010",
						 "100001100011101111010110",
						 "100001100011101011011010",
						 "100001100011100111011110",
						 "100001100011100011100010",
						 "100001100011011111100110",
						 "100001100011011011101010",
						 "100001100011010111101110",
						 "100001100011010011110010",
						 "100001100001101011111000",
						 "100001100001100111111100",
						 "100001100001100100000000",
						 "100001100001100000000100",
						 "100001100001011100001000",
						 "100001100001011000001100",
						 "100001100001010100010000",
						 "100001100001010000010100",
						 "100001100001001100011000",
						 "100001100001001000011100",
						 "100001100001000100100000",
						 "100001100001000000100100",
						 "100001100000111100101000",
						 "100001100000111000101100",
						 "100001100000110100110000",
						 "100001100000110000110100",
						 "100001100001101011111000",
						 "100001100001100111111100",
						 "100001100001100100000000",
						 "100001100001100000000100",
						 "100001100001011100001000",
						 "100001100001011000001100",
						 "100001100001010100010000",
						 "100001100001010000010100",
						 "100001100001001100011000",
						 "100001100001001000011100",
						 "100001100001000100100000",
						 "100001100001000000100100",
						 "100001100000111100101000",
						 "100001100000111000101100",
						 "100001100000110100110000",
						 "100001100000110000110100",
						 "100001011111001000111010",
						 "100001011111000100111110",
						 "100001011111000001000010",
						 "100001011110111101000110",
						 "100001011110111001001010",
						 "100001011110110101001110",
						 "100001011110110001010010",
						 "100001011110101101010110",
						 "100001011110101001011010",
						 "100001011110100101011110",
						 "100001011110100001100010",
						 "100001011110011101100110",
						 "100001011110011001101010",
						 "100001011110010101101110",
						 "100001011110010001110010",
						 "100001011110001101110110",
						 "100001011111001000111010",
						 "100001011111000100111110",
						 "100001011111000001000010",
						 "100001011110111101000110",
						 "100001011110111001001010",
						 "100001011110110101001110",
						 "100001011110110001010010",
						 "100001011110101101010110",
						 "100001011110101001011010",
						 "100001011110100101011110",
						 "100001011110100001100010",
						 "100001011110011101100110",
						 "100001011110011001101010",
						 "100001011110010101101110",
						 "100001011110010001110010",
						 "100001011110001101110110",
						 "100001011111001000111010",
						 "100001011111000100111110",
						 "100001011111000001000010",
						 "100001011110111101000110",
						 "100001011110111001001010",
						 "100001011110110101001110",
						 "100001011110110001010010",
						 "100001011110101101010110",
						 "100001011110101001011010",
						 "100001011110100101011110",
						 "100001011110100001100010",
						 "100001011110011101100110",
						 "100001011110011001101010",
						 "100001011110010101101110",
						 "100001011110010001110010",
						 "100001011110001101110110",
						 "100001011100100101111100",
						 "100001011100100010000000",
						 "100001011100011110000100",
						 "100001011100011010001000",
						 "100001011100010110001100",
						 "100001011100010010010000",
						 "100001011100001110010100",
						 "100001011100001010011000",
						 "100001011100000110011100",
						 "100001011100000010100000",
						 "100001011011111110100100",
						 "100001011011111010101000",
						 "100001011011110110101100",
						 "100001011011110010110000",
						 "100001011011101110110100",
						 "100001011011101010111000",
						 "100001011100100101111100",
						 "100001011100100010000000",
						 "100001011100011110000100",
						 "100001011100011010001000",
						 "100001011100010110001100",
						 "100001011100010010010000",
						 "100001011100001110010100",
						 "100001011100001010011000",
						 "100001011100000110011100",
						 "100001011100000010100000",
						 "100001011011111110100100",
						 "100001011011111010101000",
						 "100001011011110110101100",
						 "100001011011110010110000",
						 "100001011011101110110100",
						 "100001011011101010111000",
						 "100001011010000010111110",
						 "100001011001111111000010",
						 "100001011001111011000110",
						 "100001011001110111001010",
						 "100001011001110011001110",
						 "100001011001101111010010",
						 "100001011001101011010110",
						 "100001011001100111011010",
						 "100001011001100011011110",
						 "100001011001011111100010",
						 "100001011001011011100110",
						 "100001011001010111101010",
						 "100001011001010011101110",
						 "100001011001001111110010",
						 "100001011001001011110110",
						 "100001011001000111111010",
						 "100001011010000011001101",
						 "100001011001111111010000",
						 "100001011001111011010011",
						 "100001011001110111010110",
						 "100001011001110011011001",
						 "100001011001101111011100",
						 "100001011001101011011111",
						 "100001011001100111100010",
						 "100001011001100011100101",
						 "100001011001011111101000",
						 "100001011001011011101011",
						 "100001011001010111101110",
						 "100001011001010011110001",
						 "100001011001001111110100",
						 "100001011001001011110111",
						 "100001011001000111111010",
						 "100001011010000011001101",
						 "100001011001111111010000",
						 "100001011001111011010011",
						 "100001011001110111010110",
						 "100001011001110011011001",
						 "100001011001101111011100",
						 "100001011001101011011111",
						 "100001011001100111100010",
						 "100001011001100011100101",
						 "100001011001011111101000",
						 "100001011001011011101011",
						 "100001011001010111101110",
						 "100001011001010011110001",
						 "100001011001001111110100",
						 "100001011001001011110111",
						 "100001011001000111111010",
						 "100001010111100000001111",
						 "100001010111011100010010",
						 "100001010111011000010101",
						 "100001010111010100011000",
						 "100001010111010000011011",
						 "100001010111001100011110",
						 "100001010111001000100001",
						 "100001010111000100100100",
						 "100001010111000000100111",
						 "100001010110111100101010",
						 "100001010110111000101101",
						 "100001010110110100110000",
						 "100001010110110000110011",
						 "100001010110101100110110",
						 "100001010110101000111001",
						 "100001010110100100111100",
						 "100001010111100000001111",
						 "100001010111011100010010",
						 "100001010111011000010101",
						 "100001010111010100011000",
						 "100001010111010000011011",
						 "100001010111001100011110",
						 "100001010111001000100001",
						 "100001010111000100100100",
						 "100001010111000000100111",
						 "100001010110111100101010",
						 "100001010110111000101101",
						 "100001010110110100110000",
						 "100001010110110000110011",
						 "100001010110101100110110",
						 "100001010110101000111001",
						 "100001010110100100111100",
						 "100001010111100000001111",
						 "100001010111011100010010",
						 "100001010111011000010101",
						 "100001010111010100011000",
						 "100001010111010000011011",
						 "100001010111001100011110",
						 "100001010111001000100001",
						 "100001010111000100100100",
						 "100001010111000000100111",
						 "100001010110111100101010",
						 "100001010110111000101101",
						 "100001010110110100110000",
						 "100001010110110000110011",
						 "100001010110101100110110",
						 "100001010110101000111001",
						 "100001010110100100111100",
						 "100001010100111101010001",
						 "100001010100111001010100",
						 "100001010100110101010111",
						 "100001010100110001011010",
						 "100001010100101101011101",
						 "100001010100101001100000",
						 "100001010100100101100011",
						 "100001010100100001100110",
						 "100001010100011101101001",
						 "100001010100011001101100",
						 "100001010100010101101111",
						 "100001010100010001110010",
						 "100001010100001101110101",
						 "100001010100001001111000",
						 "100001010100000101111011",
						 "100001010100000001111110",
						 "100001010100111101010001",
						 "100001010100111001010100",
						 "100001010100110101010111",
						 "100001010100110001011010",
						 "100001010100101101011101",
						 "100001010100101001100000",
						 "100001010100100101100011",
						 "100001010100100001100110",
						 "100001010100011101101001",
						 "100001010100011001101100",
						 "100001010100010101101111",
						 "100001010100010001110010",
						 "100001010100001101110101",
						 "100001010100001001111000",
						 "100001010100000101111011",
						 "100001010100000001111110",
						 "100001010010011010010011",
						 "100001010010010110010110",
						 "100001010010010010011001",
						 "100001010010001110011100",
						 "100001010010001010011111",
						 "100001010010000110100010",
						 "100001010010000010100101",
						 "100001010001111110101000",
						 "100001010001111010101011",
						 "100001010001110110101110",
						 "100001010001110010110001",
						 "100001010001101110110100",
						 "100001010001101010110111",
						 "100001010001100110111010",
						 "100001010001100010111101",
						 "100001010001011111000000",
						 "100001010010011010010011",
						 "100001010010010110010110",
						 "100001010010010010011001",
						 "100001010010001110011100",
						 "100001010010001010011111",
						 "100001010010000110100010",
						 "100001010010000010100101",
						 "100001010001111110101000",
						 "100001010001111010101011",
						 "100001010001110110101110",
						 "100001010001110010110001",
						 "100001010001101110110100",
						 "100001010001101010110111",
						 "100001010001100110111010",
						 "100001010001100010111101",
						 "100001010001011111000000",
						 "100001010010011010010011",
						 "100001010010010110010110",
						 "100001010010010010011001",
						 "100001010010001110011100",
						 "100001010010001010011111",
						 "100001010010000110100010",
						 "100001010010000010100101",
						 "100001010001111110101000",
						 "100001010001111010101011",
						 "100001010001110110101110",
						 "100001010001110010110001",
						 "100001010001101110110100",
						 "100001010001101010110111",
						 "100001010001100110111010",
						 "100001010001100010111101",
						 "100001010001011111000000",
						 "100001001111110111010101",
						 "100001001111110011011000",
						 "100001001111101111011011",
						 "100001001111101011011110",
						 "100001001111100111100001",
						 "100001001111100011100100",
						 "100001001111011111100111",
						 "100001001111011011101010",
						 "100001001111010111101101",
						 "100001001111010011110000",
						 "100001001111001111110011",
						 "100001001111001011110110",
						 "100001001111000111111001",
						 "100001001111000011111100",
						 "100001001110111111111111",
						 "100001001110111100000010",
						 "100001001111110111010101",
						 "100001001111110011011000",
						 "100001001111101111011011",
						 "100001001111101011011110",
						 "100001001111100111100001",
						 "100001001111100011100100",
						 "100001001111011111100111",
						 "100001001111011011101010",
						 "100001001111010111101101",
						 "100001001111010011110000",
						 "100001001111001111110011",
						 "100001001111001011110110",
						 "100001001111000111111001",
						 "100001001111000011111100",
						 "100001001110111111111111",
						 "100001001110111100000010",
						 "100001001101010100010111",
						 "100001001101010000011010",
						 "100001001101001100011101",
						 "100001001101001000100000",
						 "100001001101000100100011",
						 "100001001101000000100110",
						 "100001001100111100101001",
						 "100001001100111000101100",
						 "100001001100110100101111",
						 "100001001100110000110010",
						 "100001001100101100110101",
						 "100001001100101000111000",
						 "100001001100100100111011",
						 "100001001100100000111110",
						 "100001001100011101000001",
						 "100001001100011001000100",
						 "100001001101010100010111",
						 "100001001101010000011010",
						 "100001001101001100011101",
						 "100001001101001000100000",
						 "100001001101000100100011",
						 "100001001101000000100110",
						 "100001001100111100101001",
						 "100001001100111000101100",
						 "100001001100110100101111",
						 "100001001100110000110010",
						 "100001001100101100110101",
						 "100001001100101000111000",
						 "100001001100100100111011",
						 "100001001100100000111110",
						 "100001001100011101000001",
						 "100001001100011001000100",
						 "100001001101010100010111",
						 "100001001101010000011010",
						 "100001001101001100011101",
						 "100001001101001000100000",
						 "100001001101000100100011",
						 "100001001101000000100110",
						 "100001001100111100101001",
						 "100001001100111000101100",
						 "100001001100110100101111",
						 "100001001100110000110010",
						 "100001001100101100110101",
						 "100001001100101000111000",
						 "100001001100100100111011",
						 "100001001100100000111110",
						 "100001001100011101000001",
						 "100001001100011001000100",
						 "100001001010110001011001",
						 "100001001010101101011100",
						 "100001001010101001011111",
						 "100001001010100101100010",
						 "100001001010100001100101",
						 "100001001010011101101000",
						 "100001001010011001101011",
						 "100001001010010101101110",
						 "100001001010010001110001",
						 "100001001010001101110100",
						 "100001001010001001110111",
						 "100001001010000101111010",
						 "100001001010000001111101",
						 "100001001001111110000000",
						 "100001001001111010000011",
						 "100001001001110110000110",
						 "100001001010110001011001",
						 "100001001010101101011100",
						 "100001001010101001011111",
						 "100001001010100101100010",
						 "100001001010100001100101",
						 "100001001010011101101000",
						 "100001001010011001101011",
						 "100001001010010101101110",
						 "100001001010010001110001",
						 "100001001010001101110100",
						 "100001001010001001110111",
						 "100001001010000101111010",
						 "100001001010000001111101",
						 "100001001001111110000000",
						 "100001001001111010000011",
						 "100001001001110110000110",
						 "100001001000001110011011",
						 "100001001000001010011110",
						 "100001001000000110100001",
						 "100001001000000010100100",
						 "100001000111111110100111",
						 "100001000111111010101010",
						 "100001000111110110101101",
						 "100001000111110010110000",
						 "100001000111101110110011",
						 "100001000111101010110110",
						 "100001000111100110111001",
						 "100001000111100010111100",
						 "100001000111011110111111",
						 "100001000111011011000010",
						 "100001000111010111000101",
						 "100001000111010011001000",
						 "100001001000001110011011",
						 "100001001000001010011110",
						 "100001001000000110100001",
						 "100001001000000010100100",
						 "100001000111111110100111",
						 "100001000111111010101010",
						 "100001000111110110101101",
						 "100001000111110010110000",
						 "100001000111101110110011",
						 "100001000111101010110110",
						 "100001000111100110111001",
						 "100001000111100010111100",
						 "100001000111011110111111",
						 "100001000111011011000010",
						 "100001000111010111000101",
						 "100001000111010011001000",
						 "100001001000001110011011",
						 "100001001000001010011110",
						 "100001001000000110100001",
						 "100001001000000010100100",
						 "100001000111111110100111",
						 "100001000111111010101010",
						 "100001000111110110101101",
						 "100001000111110010110000",
						 "100001000111101110110011",
						 "100001000111101010110110",
						 "100001000111100110111001",
						 "100001000111100010111100",
						 "100001000111011110111111",
						 "100001000111011011000010",
						 "100001000111010111000101",
						 "100001000111010011001000",
						 "100001000101101011101100",
						 "100001000101100111101110",
						 "100001000101100011110000",
						 "100001000101011111110010",
						 "100001000101011011110100",
						 "100001000101010111110110",
						 "100001000101010011111000",
						 "100001000101001111111010",
						 "100001000101001011111100",
						 "100001000101000111111110",
						 "100001000101000100000000",
						 "100001000101000000000010",
						 "100001000100111100000100",
						 "100001000100111000000110",
						 "100001000100110100001000",
						 "100001000100110000001010",
						 "100001000101101011101100",
						 "100001000101100111101110",
						 "100001000101100011110000",
						 "100001000101011111110010",
						 "100001000101011011110100",
						 "100001000101010111110110",
						 "100001000101010011111000",
						 "100001000101001111111010",
						 "100001000101001011111100",
						 "100001000101000111111110",
						 "100001000101000100000000",
						 "100001000101000000000010",
						 "100001000100111100000100",
						 "100001000100111000000110",
						 "100001000100110100001000",
						 "100001000100110000001010",
						 "100001000101101011101100",
						 "100001000101100111101110",
						 "100001000101100011110000",
						 "100001000101011111110010",
						 "100001000101011011110100",
						 "100001000101010111110110",
						 "100001000101010011111000",
						 "100001000101001111111010",
						 "100001000101001011111100",
						 "100001000101000111111110",
						 "100001000101000100000000",
						 "100001000101000000000010",
						 "100001000100111100000100",
						 "100001000100111000000110",
						 "100001000100110100001000",
						 "100001000100110000001010",
						 "100001000011001000101110",
						 "100001000011000100110000",
						 "100001000011000000110010",
						 "100001000010111100110100",
						 "100001000010111000110110",
						 "100001000010110100111000",
						 "100001000010110000111010",
						 "100001000010101100111100",
						 "100001000010101000111110",
						 "100001000010100101000000",
						 "100001000010100001000010",
						 "100001000010011101000100",
						 "100001000010011001000110",
						 "100001000010010101001000",
						 "100001000010010001001010",
						 "100001000010001101001100",
						 "100001000011001000101110",
						 "100001000011000100110000",
						 "100001000011000000110010",
						 "100001000010111100110100",
						 "100001000010111000110110",
						 "100001000010110100111000",
						 "100001000010110000111010",
						 "100001000010101100111100",
						 "100001000010101000111110",
						 "100001000010100101000000",
						 "100001000010100001000010",
						 "100001000010011101000100",
						 "100001000010011001000110",
						 "100001000010010101001000",
						 "100001000010010001001010",
						 "100001000010001101001100",
						 "100001000000100101110000",
						 "100001000000100001110010",
						 "100001000000011101110100",
						 "100001000000011001110110",
						 "100001000000010101111000",
						 "100001000000010001111010",
						 "100001000000001101111100",
						 "100001000000001001111110",
						 "100001000000000110000000",
						 "100001000000000010000010",
						 "100000111111111110000100",
						 "100000111111111010000110",
						 "100000111111110110001000",
						 "100000111111110010001010",
						 "100000111111101110001100",
						 "100000111111101010001110",
						 "100001000000100101110000",
						 "100001000000100001110010",
						 "100001000000011101110100",
						 "100001000000011001110110",
						 "100001000000010101111000",
						 "100001000000010001111010",
						 "100001000000001101111100",
						 "100001000000001001111110",
						 "100001000000000110000000",
						 "100001000000000010000010",
						 "100000111111111110000100",
						 "100000111111111010000110",
						 "100000111111110110001000",
						 "100000111111110010001010",
						 "100000111111101110001100",
						 "100000111111101010001110",
						 "100001000000100101110000",
						 "100001000000100001110010",
						 "100001000000011101110100",
						 "100001000000011001110110",
						 "100001000000010101111000",
						 "100001000000010001111010",
						 "100001000000001101111100",
						 "100001000000001001111110",
						 "100001000000000110000000",
						 "100001000000000010000010",
						 "100000111111111110000100",
						 "100000111111111010000110",
						 "100000111111110110001000",
						 "100000111111110010001010",
						 "100000111111101110001100",
						 "100000111111101010001110",
						 "100000111110000010110010",
						 "100000111101111110110100",
						 "100000111101111010110110",
						 "100000111101110110111000",
						 "100000111101110010111010",
						 "100000111101101110111100",
						 "100000111101101010111110",
						 "100000111101100111000000",
						 "100000111101100011000010",
						 "100000111101011111000100",
						 "100000111101011011000110",
						 "100000111101010111001000",
						 "100000111101010011001010",
						 "100000111101001111001100",
						 "100000111101001011001110",
						 "100000111101000111010000",
						 "100000111110000010110010",
						 "100000111101111110110100",
						 "100000111101111010110110",
						 "100000111101110110111000",
						 "100000111101110010111010",
						 "100000111101101110111100",
						 "100000111101101010111110",
						 "100000111101100111000000",
						 "100000111101100011000010",
						 "100000111101011111000100",
						 "100000111101011011000110",
						 "100000111101010111001000",
						 "100000111101010011001010",
						 "100000111101001111001100",
						 "100000111101001011001110",
						 "100000111101000111010000",
						 "100000111011011111110100",
						 "100000111011011011110110",
						 "100000111011010111111000",
						 "100000111011010011111010",
						 "100000111011001111111100",
						 "100000111011001011111110",
						 "100000111011001000000000",
						 "100000111011000100000010",
						 "100000111011000000000100",
						 "100000111010111100000110",
						 "100000111010111000001000",
						 "100000111010110100001010",
						 "100000111010110000001100",
						 "100000111010101100001110",
						 "100000111010101000010000",
						 "100000111010100100010010",
						 "100000111011011111110100",
						 "100000111011011011110110",
						 "100000111011010111111000",
						 "100000111011010011111010",
						 "100000111011001111111100",
						 "100000111011001011111110",
						 "100000111011001000000000",
						 "100000111011000100000010",
						 "100000111011000000000100",
						 "100000111010111100000110",
						 "100000111010111000001000",
						 "100000111010110100001010",
						 "100000111010110000001100",
						 "100000111010101100001110",
						 "100000111010101000010000",
						 "100000111010100100010010",
						 "100000111011011111110100",
						 "100000111011011011110110",
						 "100000111011010111111000",
						 "100000111011010011111010",
						 "100000111011001111111100",
						 "100000111011001011111110",
						 "100000111011001000000000",
						 "100000111011000100000010",
						 "100000111011000000000100",
						 "100000111010111100000110",
						 "100000111010111000001000",
						 "100000111010110100001010",
						 "100000111010110000001100",
						 "100000111010101100001110",
						 "100000111010101000010000",
						 "100000111010100100010010",
						 "100000111000111100110110",
						 "100000111000111000111000",
						 "100000111000110100111010",
						 "100000111000110000111100",
						 "100000111000101100111110",
						 "100000111000101001000000",
						 "100000111000100101000010",
						 "100000111000100001000100",
						 "100000111000011101000110",
						 "100000111000011001001000",
						 "100000111000010101001010",
						 "100000111000010001001100",
						 "100000111000001101001110",
						 "100000111000001001010000",
						 "100000111000000101010010",
						 "100000111000000001010100",
						 "100000111000111100110110",
						 "100000111000111000111000",
						 "100000111000110100111010",
						 "100000111000110000111100",
						 "100000111000101100111110",
						 "100000111000101001000000",
						 "100000111000100101000010",
						 "100000111000100001000100",
						 "100000111000011101000110",
						 "100000111000011001001000",
						 "100000111000010101001010",
						 "100000111000010001001100",
						 "100000111000001101001110",
						 "100000111000001001010000",
						 "100000111000000101010010",
						 "100000111000000001010100",
						 "100000110110011001111000",
						 "100000110110010101111010",
						 "100000110110010001111100",
						 "100000110110001101111110",
						 "100000110110001010000000",
						 "100000110110000110000010",
						 "100000110110000010000100",
						 "100000110101111110000110",
						 "100000110101111010001000",
						 "100000110101110110001010",
						 "100000110101110010001100",
						 "100000110101101110001110",
						 "100000110101101010010000",
						 "100000110101100110010010",
						 "100000110101100010010100",
						 "100000110101011110010110",
						 "100000110110011001111000",
						 "100000110110010101111010",
						 "100000110110010001111100",
						 "100000110110001101111110",
						 "100000110110001010000000",
						 "100000110110000110000010",
						 "100000110110000010000100",
						 "100000110101111110000110",
						 "100000110101111010001000",
						 "100000110101110110001010",
						 "100000110101110010001100",
						 "100000110101101110001110",
						 "100000110101101010010000",
						 "100000110101100110010010",
						 "100000110101100010010100",
						 "100000110101011110010110",
						 "100000110110011001111000",
						 "100000110110010101111010",
						 "100000110110010001111100",
						 "100000110110001101111110",
						 "100000110110001010000000",
						 "100000110110000110000010",
						 "100000110110000010000100",
						 "100000110101111110000110",
						 "100000110101111010001000",
						 "100000110101110110001010",
						 "100000110101110010001100",
						 "100000110101101110001110",
						 "100000110101101010010000",
						 "100000110101100110010010",
						 "100000110101100010010100",
						 "100000110101011110010110",
						 "100000110011110110111010",
						 "100000110011110010111100",
						 "100000110011101110111110",
						 "100000110011101011000000",
						 "100000110011100111000010",
						 "100000110011100011000100",
						 "100000110011011111000110",
						 "100000110011011011001000",
						 "100000110011010111001010",
						 "100000110011010011001100",
						 "100000110011001111001110",
						 "100000110011001011010000",
						 "100000110011000111010010",
						 "100000110011000011010100",
						 "100000110010111111010110",
						 "100000110010111011011000",
						 "100000110011110110111010",
						 "100000110011110010111100",
						 "100000110011101110111110",
						 "100000110011101011000000",
						 "100000110011100111000010",
						 "100000110011100011000100",
						 "100000110011011111000110",
						 "100000110011011011001000",
						 "100000110011010111001010",
						 "100000110011010011001100",
						 "100000110011001111001110",
						 "100000110011001011010000",
						 "100000110011000111010010",
						 "100000110011000011010100",
						 "100000110010111111010110",
						 "100000110010111011011000",
						 "100000110011110110111010",
						 "100000110011110010111100",
						 "100000110011101110111110",
						 "100000110011101011000000",
						 "100000110011100111000010",
						 "100000110011100011000100",
						 "100000110011011111000110",
						 "100000110011011011001000",
						 "100000110011010111001010",
						 "100000110011010011001100",
						 "100000110011001111001110",
						 "100000110011001011010000",
						 "100000110011000111010010",
						 "100000110011000011010100",
						 "100000110010111111010110",
						 "100000110010111011011000",
						 "100000110001010011111100",
						 "100000110001001111111110",
						 "100000110001001100000000",
						 "100000110001001000000010",
						 "100000110001000100000100",
						 "100000110001000000000110",
						 "100000110000111100001000",
						 "100000110000111000001010",
						 "100000110000110100001100",
						 "100000110000110000001110",
						 "100000110000101100010000",
						 "100000110000101000010010",
						 "100000110000100100010100",
						 "100000110000100000010110",
						 "100000110000011100011000",
						 "100000110000011000011010",
						 "100000110001010011111100",
						 "100000110001001111111110",
						 "100000110001001100000000",
						 "100000110001001000000010",
						 "100000110001000100000100",
						 "100000110001000000000110",
						 "100000110000111100001000",
						 "100000110000111000001010",
						 "100000110000110100001100",
						 "100000110000110000001110",
						 "100000110000101100010000",
						 "100000110000101000010010",
						 "100000110000100100010100",
						 "100000110000100000010110",
						 "100000110000011100011000",
						 "100000110000011000011010",
						 "100000101110110000111110",
						 "100000101110101101000000",
						 "100000101110101001000010",
						 "100000101110100101000100",
						 "100000101110100001000110",
						 "100000101110011101001000",
						 "100000101110011001001010",
						 "100000101110010101001100",
						 "100000101110010001001110",
						 "100000101110001101010000",
						 "100000101110001001010010",
						 "100000101110000101010100",
						 "100000101110000001010110",
						 "100000101101111101011000",
						 "100000101101111001011010",
						 "100000101101110101011100",
						 "100000101110110000111110",
						 "100000101110101101000000",
						 "100000101110101001000010",
						 "100000101110100101000100",
						 "100000101110100001000110",
						 "100000101110011101001000",
						 "100000101110011001001010",
						 "100000101110010101001100",
						 "100000101110010001001110",
						 "100000101110001101010000",
						 "100000101110001001010010",
						 "100000101110000101010100",
						 "100000101110000001010110",
						 "100000101101111101011000",
						 "100000101101111001011010",
						 "100000101101110101011100",
						 "100000101110110000111110",
						 "100000101110101101000000",
						 "100000101110101001000010",
						 "100000101110100101000100",
						 "100000101110100001000110",
						 "100000101110011101001000",
						 "100000101110011001001010",
						 "100000101110010101001100",
						 "100000101110010001001110",
						 "100000101110001101010000",
						 "100000101110001001010010",
						 "100000101110000101010100",
						 "100000101110000001010110",
						 "100000101101111101011000",
						 "100000101101111001011010",
						 "100000101101110101011100",
						 "100000101100001110000000",
						 "100000101100001010000010",
						 "100000101100000110000100",
						 "100000101100000010000110",
						 "100000101011111110001000",
						 "100000101011111010001010",
						 "100000101011110110001100",
						 "100000101011110010001110",
						 "100000101011101110010000",
						 "100000101011101010010010",
						 "100000101011100110010100",
						 "100000101011100010010110",
						 "100000101011011110011000",
						 "100000101011011010011010",
						 "100000101011010110011100",
						 "100000101011010010011110",
						 "100000101100001110000000",
						 "100000101100001010000010",
						 "100000101100000110000100",
						 "100000101100000010000110",
						 "100000101011111110001000",
						 "100000101011111010001010",
						 "100000101011110110001100",
						 "100000101011110010001110",
						 "100000101011101110010000",
						 "100000101011101010010010",
						 "100000101011100110010100",
						 "100000101011100010010110",
						 "100000101011011110011000",
						 "100000101011011010011010",
						 "100000101011010110011100",
						 "100000101011010010011110",
						 "100000101001101011000010",
						 "100000101001100111000100",
						 "100000101001100011000110",
						 "100000101001011111001000",
						 "100000101001011011001010",
						 "100000101001010111001100",
						 "100000101001010011001110",
						 "100000101001001111010000",
						 "100000101001001011010010",
						 "100000101001000111010100",
						 "100000101001000011010110",
						 "100000101000111111011000",
						 "100000101000111011011010",
						 "100000101000110111011100",
						 "100000101000110011011110",
						 "100000101000101111100000",
						 "100000101001101011000010",
						 "100000101001100111000100",
						 "100000101001100011000110",
						 "100000101001011111001000",
						 "100000101001011011001010",
						 "100000101001010111001100",
						 "100000101001010011001110",
						 "100000101001001111010000",
						 "100000101001001011010010",
						 "100000101001000111010100",
						 "100000101001000011010110",
						 "100000101000111111011000",
						 "100000101000111011011010",
						 "100000101000110111011100",
						 "100000101000110011011110",
						 "100000101000101111100000",
						 "100000101001101011010001",
						 "100000101001100111010010",
						 "100000101001100011010011",
						 "100000101001011111010100",
						 "100000101001011011010101",
						 "100000101001010111010110",
						 "100000101001010011010111",
						 "100000101001001111011000",
						 "100000101001001011011001",
						 "100000101001000111011010",
						 "100000101001000011011011",
						 "100000101000111111011100",
						 "100000101000111011011101",
						 "100000101000110111011110",
						 "100000101000110011011111",
						 "100000101000101111100000",
						 "100000100111001000010011",
						 "100000100111000100010100",
						 "100000100111000000010101",
						 "100000100110111100010110",
						 "100000100110111000010111",
						 "100000100110110100011000",
						 "100000100110110000011001",
						 "100000100110101100011010",
						 "100000100110101000011011",
						 "100000100110100100011100",
						 "100000100110100000011101",
						 "100000100110011100011110",
						 "100000100110011000011111",
						 "100000100110010100100000",
						 "100000100110010000100001",
						 "100000100110001100100010",
						 "100000100111001000010011",
						 "100000100111000100010100",
						 "100000100111000000010101",
						 "100000100110111100010110",
						 "100000100110111000010111",
						 "100000100110110100011000",
						 "100000100110110000011001",
						 "100000100110101100011010",
						 "100000100110101000011011",
						 "100000100110100100011100",
						 "100000100110100000011101",
						 "100000100110011100011110",
						 "100000100110011000011111",
						 "100000100110010100100000",
						 "100000100110010000100001",
						 "100000100110001100100010",
						 "100000100100100101010101",
						 "100000100100100001010110",
						 "100000100100011101010111",
						 "100000100100011001011000",
						 "100000100100010101011001",
						 "100000100100010001011010",
						 "100000100100001101011011",
						 "100000100100001001011100",
						 "100000100100000101011101",
						 "100000100100000001011110",
						 "100000100011111101011111",
						 "100000100011111001100000",
						 "100000100011110101100001",
						 "100000100011110001100010",
						 "100000100011101101100011",
						 "100000100011101001100100",
						 "100000100100100101010101",
						 "100000100100100001010110",
						 "100000100100011101010111",
						 "100000100100011001011000",
						 "100000100100010101011001",
						 "100000100100010001011010",
						 "100000100100001101011011",
						 "100000100100001001011100",
						 "100000100100000101011101",
						 "100000100100000001011110",
						 "100000100011111101011111",
						 "100000100011111001100000",
						 "100000100011110101100001",
						 "100000100011110001100010",
						 "100000100011101101100011",
						 "100000100011101001100100",
						 "100000100100100101010101",
						 "100000100100100001010110",
						 "100000100100011101010111",
						 "100000100100011001011000",
						 "100000100100010101011001",
						 "100000100100010001011010",
						 "100000100100001101011011",
						 "100000100100001001011100",
						 "100000100100000101011101",
						 "100000100100000001011110",
						 "100000100011111101011111",
						 "100000100011111001100000",
						 "100000100011110101100001",
						 "100000100011110001100010",
						 "100000100011101101100011",
						 "100000100011101001100100",
						 "100000100010000010010111",
						 "100000100001111110011000",
						 "100000100001111010011001",
						 "100000100001110110011010",
						 "100000100001110010011011",
						 "100000100001101110011100",
						 "100000100001101010011101",
						 "100000100001100110011110",
						 "100000100001100010011111",
						 "100000100001011110100000",
						 "100000100001011010100001",
						 "100000100001010110100010",
						 "100000100001010010100011",
						 "100000100001001110100100",
						 "100000100001001010100101",
						 "100000100001000110100110",
						 "100000100010000010010111",
						 "100000100001111110011000",
						 "100000100001111010011001",
						 "100000100001110110011010",
						 "100000100001110010011011",
						 "100000100001101110011100",
						 "100000100001101010011101",
						 "100000100001100110011110",
						 "100000100001100010011111",
						 "100000100001011110100000",
						 "100000100001011010100001",
						 "100000100001010110100010",
						 "100000100001010010100011",
						 "100000100001001110100100",
						 "100000100001001010100101",
						 "100000100001000110100110",
						 "100000100010000010010111",
						 "100000100001111110011000",
						 "100000100001111010011001",
						 "100000100001110110011010",
						 "100000100001110010011011",
						 "100000100001101110011100",
						 "100000100001101010011101",
						 "100000100001100110011110",
						 "100000100001100010011111",
						 "100000100001011110100000",
						 "100000100001011010100001",
						 "100000100001010110100010",
						 "100000100001010010100011",
						 "100000100001001110100100",
						 "100000100001001010100101",
						 "100000100001000110100110",
						 "100000011111011111011001",
						 "100000011111011011011010",
						 "100000011111010111011011",
						 "100000011111010011011100",
						 "100000011111001111011101",
						 "100000011111001011011110",
						 "100000011111000111011111",
						 "100000011111000011100000",
						 "100000011110111111100001",
						 "100000011110111011100010",
						 "100000011110110111100011",
						 "100000011110110011100100",
						 "100000011110101111100101",
						 "100000011110101011100110",
						 "100000011110100111100111",
						 "100000011110100011101000",
						 "100000011111011111011001",
						 "100000011111011011011010",
						 "100000011111010111011011",
						 "100000011111010011011100",
						 "100000011111001111011101",
						 "100000011111001011011110",
						 "100000011111000111011111",
						 "100000011111000011100000",
						 "100000011110111111100001",
						 "100000011110111011100010",
						 "100000011110110111100011",
						 "100000011110110011100100",
						 "100000011110101111100101",
						 "100000011110101011100110",
						 "100000011110100111100111",
						 "100000011110100011101000",
						 "100000011100111100011011",
						 "100000011100111000011100",
						 "100000011100110100011101",
						 "100000011100110000011110",
						 "100000011100101100011111",
						 "100000011100101000100000",
						 "100000011100100100100001",
						 "100000011100100000100010",
						 "100000011100011100100011",
						 "100000011100011000100100",
						 "100000011100010100100101",
						 "100000011100010000100110",
						 "100000011100001100100111",
						 "100000011100001000101000",
						 "100000011100000100101001",
						 "100000011100000000101010",
						 "100000011100111100011011",
						 "100000011100111000011100",
						 "100000011100110100011101",
						 "100000011100110000011110",
						 "100000011100101100011111",
						 "100000011100101000100000",
						 "100000011100100100100001",
						 "100000011100100000100010",
						 "100000011100011100100011",
						 "100000011100011000100100",
						 "100000011100010100100101",
						 "100000011100010000100110",
						 "100000011100001100100111",
						 "100000011100001000101000",
						 "100000011100000100101001",
						 "100000011100000000101010",
						 "100000011100111100011011",
						 "100000011100111000011100",
						 "100000011100110100011101",
						 "100000011100110000011110",
						 "100000011100101100011111",
						 "100000011100101000100000",
						 "100000011100100100100001",
						 "100000011100100000100010",
						 "100000011100011100100011",
						 "100000011100011000100100",
						 "100000011100010100100101",
						 "100000011100010000100110",
						 "100000011100001100100111",
						 "100000011100001000101000",
						 "100000011100000100101001",
						 "100000011100000000101010",
						 "100000011010011001011101",
						 "100000011010010101011110",
						 "100000011010010001011111",
						 "100000011010001101100000",
						 "100000011010001001100001",
						 "100000011010000101100010",
						 "100000011010000001100011",
						 "100000011001111101100100",
						 "100000011001111001100101",
						 "100000011001110101100110",
						 "100000011001110001100111",
						 "100000011001101101101000",
						 "100000011001101001101001",
						 "100000011001100101101010",
						 "100000011001100001101011",
						 "100000011001011101101100",
						 "100000011010011001011101",
						 "100000011010010101011110",
						 "100000011010010001011111",
						 "100000011010001101100000",
						 "100000011010001001100001",
						 "100000011010000101100010",
						 "100000011010000001100011",
						 "100000011001111101100100",
						 "100000011001111001100101",
						 "100000011001110101100110",
						 "100000011001110001100111",
						 "100000011001101101101000",
						 "100000011001101001101001",
						 "100000011001100101101010",
						 "100000011001100001101011",
						 "100000011001011101101100",
						 "100000010111110110011111",
						 "100000010111110010100000",
						 "100000010111101110100001",
						 "100000010111101010100010",
						 "100000010111100110100011",
						 "100000010111100010100100",
						 "100000010111011110100101",
						 "100000010111011010100110",
						 "100000010111010110100111",
						 "100000010111010010101000",
						 "100000010111001110101001",
						 "100000010111001010101010",
						 "100000010111000110101011",
						 "100000010111000010101100",
						 "100000010110111110101101",
						 "100000010110111010101110",
						 "100000010111110110011111",
						 "100000010111110010100000",
						 "100000010111101110100001",
						 "100000010111101010100010",
						 "100000010111100110100011",
						 "100000010111100010100100",
						 "100000010111011110100101",
						 "100000010111011010100110",
						 "100000010111010110100111",
						 "100000010111010010101000",
						 "100000010111001110101001",
						 "100000010111001010101010",
						 "100000010111000110101011",
						 "100000010111000010101100",
						 "100000010110111110101101",
						 "100000010110111010101110",
						 "100000010111110110011111",
						 "100000010111110010100000",
						 "100000010111101110100001",
						 "100000010111101010100010",
						 "100000010111100110100011",
						 "100000010111100010100100",
						 "100000010111011110100101",
						 "100000010111011010100110",
						 "100000010111010110100111",
						 "100000010111010010101000",
						 "100000010111001110101001",
						 "100000010111001010101010",
						 "100000010111000110101011",
						 "100000010111000010101100",
						 "100000010110111110101101",
						 "100000010110111010101110",
						 "100000010101010011100001",
						 "100000010101001111100010",
						 "100000010101001011100011",
						 "100000010101000111100100",
						 "100000010101000011100101",
						 "100000010100111111100110",
						 "100000010100111011100111",
						 "100000010100110111101000",
						 "100000010100110011101001",
						 "100000010100101111101010",
						 "100000010100101011101011",
						 "100000010100100111101100",
						 "100000010100100011101101",
						 "100000010100011111101110",
						 "100000010100011011101111",
						 "100000010100010111110000",
						 "100000010101010011100001",
						 "100000010101001111100010",
						 "100000010101001011100011",
						 "100000010101000111100100",
						 "100000010101000011100101",
						 "100000010100111111100110",
						 "100000010100111011100111",
						 "100000010100110111101000",
						 "100000010100110011101001",
						 "100000010100101111101010",
						 "100000010100101011101011",
						 "100000010100100111101100",
						 "100000010100100011101101",
						 "100000010100011111101110",
						 "100000010100011011101111",
						 "100000010100010111110000",
						 "100000010010110000100011",
						 "100000010010101100100100",
						 "100000010010101000100101",
						 "100000010010100100100110",
						 "100000010010100000100111",
						 "100000010010011100101000",
						 "100000010010011000101001",
						 "100000010010010100101010",
						 "100000010010010000101011",
						 "100000010010001100101100",
						 "100000010010001000101101",
						 "100000010010000100101110",
						 "100000010010000000101111",
						 "100000010001111100110000",
						 "100000010001111000110001",
						 "100000010001110100110010",
						 "100000010010110000100011",
						 "100000010010101100100100",
						 "100000010010101000100101",
						 "100000010010100100100110",
						 "100000010010100000100111",
						 "100000010010011100101000",
						 "100000010010011000101001",
						 "100000010010010100101010",
						 "100000010010010000101011",
						 "100000010010001100101100",
						 "100000010010001000101101",
						 "100000010010000100101110",
						 "100000010010000000101111",
						 "100000010001111100110000",
						 "100000010001111000110001",
						 "100000010001110100110010",
						 "100000010010110000100011",
						 "100000010010101100100100",
						 "100000010010101000100101",
						 "100000010010100100100110",
						 "100000010010100000100111",
						 "100000010010011100101000",
						 "100000010010011000101001",
						 "100000010010010100101010",
						 "100000010010010000101011",
						 "100000010010001100101100",
						 "100000010010001000101101",
						 "100000010010000100101110",
						 "100000010010000000101111",
						 "100000010001111100110000",
						 "100000010001111000110001",
						 "100000010001110100110010",
						 "100000010000001101100101",
						 "100000010000001001100110",
						 "100000010000000101100111",
						 "100000010000000001101000",
						 "100000001111111101101001",
						 "100000001111111001101010",
						 "100000001111110101101011",
						 "100000001111110001101100",
						 "100000001111101101101101",
						 "100000001111101001101110",
						 "100000001111100101101111",
						 "100000001111100001110000",
						 "100000001111011101110001",
						 "100000001111011001110010",
						 "100000001111010101110011",
						 "100000001111010001110100",
						 "100000010000001101100101",
						 "100000010000001001100110",
						 "100000010000000101100111",
						 "100000010000000001101000",
						 "100000001111111101101001",
						 "100000001111111001101010",
						 "100000001111110101101011",
						 "100000001111110001101100",
						 "100000001111101101101101",
						 "100000001111101001101110",
						 "100000001111100101101111",
						 "100000001111100001110000",
						 "100000001111011101110001",
						 "100000001111011001110010",
						 "100000001111010101110011",
						 "100000001111010001110100",
						 "100000001101101010100111",
						 "100000001101100110101000",
						 "100000001101100010101001",
						 "100000001101011110101010",
						 "100000001101011010101011",
						 "100000001101010110101100",
						 "100000001101010010101101",
						 "100000001101001110101110",
						 "100000001101001010101111",
						 "100000001101000110110000",
						 "100000001101000010110001",
						 "100000001100111110110010",
						 "100000001100111010110011",
						 "100000001100110110110100",
						 "100000001100110010110101",
						 "100000001100101110110110",
						 "100000001101101010100111",
						 "100000001101100110101000",
						 "100000001101100010101001",
						 "100000001101011110101010",
						 "100000001101011010101011",
						 "100000001101010110101100",
						 "100000001101010010101101",
						 "100000001101001110101110",
						 "100000001101001010101111",
						 "100000001101000110110000",
						 "100000001101000010110001",
						 "100000001100111110110010",
						 "100000001100111010110011",
						 "100000001100110110110100",
						 "100000001100110010110101",
						 "100000001100101110110110",
						 "100000001101101010100111",
						 "100000001101100110101000",
						 "100000001101100010101001",
						 "100000001101011110101010",
						 "100000001101011010101011",
						 "100000001101010110101100",
						 "100000001101010010101101",
						 "100000001101001110101110",
						 "100000001101001010101111",
						 "100000001101000110110000",
						 "100000001101000010110001",
						 "100000001100111110110010",
						 "100000001100111010110011",
						 "100000001100110110110100",
						 "100000001100110010110101",
						 "100000001100101110110110",
						 "100000001011000111101001",
						 "100000001011000011101010",
						 "100000001010111111101011",
						 "100000001010111011101100",
						 "100000001010110111101101",
						 "100000001010110011101110",
						 "100000001010101111101111",
						 "100000001010101011110000",
						 "100000001010100111110001",
						 "100000001010100011110010",
						 "100000001010011111110011",
						 "100000001010011011110100",
						 "100000001010010111110101",
						 "100000001010010011110110",
						 "100000001010001111110111",
						 "100000001010001011111000",
						 "100000001011000111101001",
						 "100000001011000011101010",
						 "100000001010111111101011",
						 "100000001010111011101100",
						 "100000001010110111101101",
						 "100000001010110011101110",
						 "100000001010101111101111",
						 "100000001010101011110000",
						 "100000001010100111110001",
						 "100000001010100011110010",
						 "100000001010011111110011",
						 "100000001010011011110100",
						 "100000001010010111110101",
						 "100000001010010011110110",
						 "100000001010001111110111",
						 "100000001010001011111000",
						 "100000001011000111101001",
						 "100000001011000011101010",
						 "100000001010111111101011",
						 "100000001010111011101100",
						 "100000001010110111101101",
						 "100000001010110011101110",
						 "100000001010101111101111",
						 "100000001010101011110000",
						 "100000001010100111110001",
						 "100000001010100011110010",
						 "100000001010011111110011",
						 "100000001010011011110100",
						 "100000001010010111110101",
						 "100000001010010011110110",
						 "100000001010001111110111",
						 "100000001010001011111000",
						 "100000001000100100101011",
						 "100000001000100000101100",
						 "100000001000011100101101",
						 "100000001000011000101110",
						 "100000001000010100101111",
						 "100000001000010000110000",
						 "100000001000001100110001",
						 "100000001000001000110010",
						 "100000001000000100110011",
						 "100000001000000000110100",
						 "100000000111111100110101",
						 "100000000111111000110110",
						 "100000000111110100110111",
						 "100000000111110000111000",
						 "100000000111101100111001",
						 "100000000111101000111010",
						 "100000001000100100101011",
						 "100000001000100000101100",
						 "100000001000011100101101",
						 "100000001000011000101110",
						 "100000001000010100101111",
						 "100000001000010000110000",
						 "100000001000001100110001",
						 "100000001000001000110010",
						 "100000001000000100110011",
						 "100000001000000000110100",
						 "100000000111111100110101",
						 "100000000111111000110110",
						 "100000000111110100110111",
						 "100000000111110000111000",
						 "100000000111101100111001",
						 "100000000111101000111010",
						 "100000000110000001101101",
						 "100000000101111101101110",
						 "100000000101111001101111",
						 "100000000101110101110000",
						 "100000000101110001110001",
						 "100000000101101101110010",
						 "100000000101101001110011",
						 "100000000101100101110100",
						 "100000000101100001110101",
						 "100000000101011101110110",
						 "100000000101011001110111",
						 "100000000101010101111000",
						 "100000000101010001111001",
						 "100000000101001101111010",
						 "100000000101001001111011",
						 "100000000101000101111100",
						 "100000000110000001101101",
						 "100000000101111101101110",
						 "100000000101111001101111",
						 "100000000101110101110000",
						 "100000000101110001110001",
						 "100000000101101101110010",
						 "100000000101101001110011",
						 "100000000101100101110100",
						 "100000000101100001110101",
						 "100000000101011101110110",
						 "100000000101011001110111",
						 "100000000101010101111000",
						 "100000000101010001111001",
						 "100000000101001101111010",
						 "100000000101001001111011",
						 "100000000101000101111100",
						 "100000000110000001101101",
						 "100000000101111101101110",
						 "100000000101111001101111",
						 "100000000101110101110000",
						 "100000000101110001110001",
						 "100000000101101101110010",
						 "100000000101101001110011",
						 "100000000101100101110100",
						 "100000000101100001110101",
						 "100000000101011101110110",
						 "100000000101011001110111",
						 "100000000101010101111000",
						 "100000000101010001111001",
						 "100000000101001101111010",
						 "100000000101001001111011",
						 "100000000101000101111100",
						 "100000000011011110101111",
						 "100000000011011010110000",
						 "100000000011010110110001",
						 "100000000011010010110010",
						 "100000000011001110110011",
						 "100000000011001010110100",
						 "100000000011000110110101",
						 "100000000011000010110110",
						 "100000000010111110110111",
						 "100000000010111010111000",
						 "100000000010110110111001",
						 "100000000010110010111010",
						 "100000000010101110111011",
						 "100000000010101010111100",
						 "100000000010100110111101",
						 "100000000010100010111110",
						 "100000000011011110101111",
						 "100000000011011010110000",
						 "100000000011010110110001",
						 "100000000011010010110010",
						 "100000000011001110110011",
						 "100000000011001010110100",
						 "100000000011000110110101",
						 "100000000011000010110110",
						 "100000000010111110110111",
						 "100000000010111010111000",
						 "100000000010110110111001",
						 "100000000010110010111010",
						 "100000000010101110111011",
						 "100000000010101010111100",
						 "100000000010100110111101",
						 "100000000010100010111110",
						 "100000000000111011110001",
						 "100000000000110111110010",
						 "100000000000110011110011",
						 "100000000000101111110100",
						 "100000000000101011110101",
						 "100000000000100111110110",
						 "100000000000100011110111",
						 "100000000000011111111000",
						 "100000000000011011111001",
						 "100000000000010111111010",
						 "100000000000010011111011",
						 "100000000000001111111100",
						 "100000000000001011111101",
						 "100000000000000111111110",
						 "100000000000000011111111",
						 "100000000000000000000000",
						 "100000000000111011110001",
						 "100000000000110111110010",
						 "100000000000110011110011",
						 "100000000000101111110100",
						 "100000000000101011110101",
						 "100000000000100111110110",
						 "100000000000100011110111",
						 "100000000000011111111000",
						 "100000000000011011111001",
						 "100000000000010111111010",
						 "100000000000010011111011",
						 "100000000000001111111100",
						 "100000000000001011111101",
						 "100000000000000111111110",
						 "100000000000000011111111",
						 "100000000000000000000000");


begin

    rom_proc: process(reset, clock)
    begin
        if reset = '1' then
            data <= (others => '0');
        elsif rising_edge(clock) then
            data <= rom(to_integer(unsigned(address)));
        end if;
    end process;

end Behaviour;